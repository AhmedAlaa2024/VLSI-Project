
// 	Sat Dec 24 03:56:12 2022
//	vlsi
//	localhost.localdomain

module register__parameterized0 (DATA_IN, DATA_OUT, clk, reset);

output [63:0] DATA_OUT;
input [63:0] DATA_IN;
input clk;
input reset;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;


AND2_X2 i_0_63 (.ZN (n_63), .A1 (reset), .A2 (DATA_IN[63]));
AND2_X1 i_0_62 (.ZN (n_62), .A1 (reset), .A2 (DATA_IN[62]));
AND2_X2 i_0_61 (.ZN (n_61), .A1 (reset), .A2 (DATA_IN[61]));
AND2_X1 i_0_60 (.ZN (n_60), .A1 (reset), .A2 (DATA_IN[60]));
AND2_X1 i_0_59 (.ZN (n_59), .A1 (reset), .A2 (DATA_IN[59]));
AND2_X2 i_0_58 (.ZN (n_58), .A1 (reset), .A2 (DATA_IN[58]));
AND2_X1 i_0_57 (.ZN (n_57), .A1 (reset), .A2 (DATA_IN[57]));
AND2_X2 i_0_56 (.ZN (n_56), .A1 (reset), .A2 (DATA_IN[56]));
AND2_X2 i_0_55 (.ZN (n_55), .A1 (reset), .A2 (DATA_IN[55]));
AND2_X2 i_0_54 (.ZN (n_54), .A1 (reset), .A2 (DATA_IN[54]));
AND2_X1 i_0_53 (.ZN (n_53), .A1 (reset), .A2 (DATA_IN[53]));
AND2_X2 i_0_52 (.ZN (n_52), .A1 (reset), .A2 (DATA_IN[52]));
AND2_X1 i_0_51 (.ZN (n_51), .A1 (reset), .A2 (DATA_IN[51]));
AND2_X1 i_0_50 (.ZN (n_50), .A1 (reset), .A2 (DATA_IN[50]));
AND2_X1 i_0_49 (.ZN (n_49), .A1 (reset), .A2 (DATA_IN[49]));
AND2_X1 i_0_48 (.ZN (n_48), .A1 (reset), .A2 (DATA_IN[48]));
AND2_X1 i_0_47 (.ZN (n_47), .A1 (reset), .A2 (DATA_IN[47]));
AND2_X1 i_0_46 (.ZN (n_46), .A1 (reset), .A2 (DATA_IN[46]));
AND2_X1 i_0_45 (.ZN (n_45), .A1 (reset), .A2 (DATA_IN[45]));
AND2_X1 i_0_44 (.ZN (n_44), .A1 (reset), .A2 (DATA_IN[44]));
AND2_X1 i_0_43 (.ZN (n_43), .A1 (reset), .A2 (DATA_IN[43]));
AND2_X1 i_0_42 (.ZN (n_42), .A1 (reset), .A2 (DATA_IN[42]));
AND2_X1 i_0_41 (.ZN (n_41), .A1 (reset), .A2 (DATA_IN[41]));
AND2_X1 i_0_40 (.ZN (n_40), .A1 (reset), .A2 (DATA_IN[40]));
AND2_X1 i_0_39 (.ZN (n_39), .A1 (reset), .A2 (DATA_IN[39]));
AND2_X1 i_0_38 (.ZN (n_38), .A1 (reset), .A2 (DATA_IN[38]));
AND2_X1 i_0_37 (.ZN (n_37), .A1 (reset), .A2 (DATA_IN[37]));
AND2_X1 i_0_36 (.ZN (n_36), .A1 (reset), .A2 (DATA_IN[36]));
AND2_X1 i_0_35 (.ZN (n_35), .A1 (reset), .A2 (DATA_IN[35]));
AND2_X1 i_0_34 (.ZN (n_34), .A1 (reset), .A2 (DATA_IN[34]));
AND2_X1 i_0_33 (.ZN (n_33), .A1 (reset), .A2 (DATA_IN[33]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (reset), .A2 (DATA_IN[32]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (reset), .A2 (DATA_IN[31]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (reset), .A2 (DATA_IN[30]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (reset), .A2 (DATA_IN[29]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (reset), .A2 (DATA_IN[28]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (reset), .A2 (DATA_IN[27]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (reset), .A2 (DATA_IN[26]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (reset), .A2 (DATA_IN[25]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (reset), .A2 (DATA_IN[24]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (reset), .A2 (DATA_IN[23]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (reset), .A2 (DATA_IN[22]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (reset), .A2 (DATA_IN[21]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (reset), .A2 (DATA_IN[20]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (reset), .A2 (DATA_IN[19]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (reset), .A2 (DATA_IN[18]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (reset), .A2 (DATA_IN[17]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (reset), .A2 (DATA_IN[16]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (reset), .A2 (DATA_IN[15]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (reset), .A2 (DATA_IN[14]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (reset), .A2 (DATA_IN[13]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (reset), .A2 (DATA_IN[12]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (reset), .A2 (DATA_IN[11]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (reset), .A2 (DATA_IN[10]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (reset), .A2 (DATA_IN[9]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (reset), .A2 (DATA_IN[8]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (reset), .A2 (DATA_IN[7]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (reset), .A2 (DATA_IN[6]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (reset), .A2 (DATA_IN[5]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (reset), .A2 (DATA_IN[4]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (reset), .A2 (DATA_IN[3]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (reset), .A2 (DATA_IN[2]));
AND2_X1 i_0_1 (.ZN (n_1), .A1 (reset), .A2 (DATA_IN[1]));
AND2_X1 i_0_0 (.ZN (n_0), .A1 (DATA_IN[0]), .A2 (reset));
DFF_X1 \DATA_reg[0]  (.Q (DATA_OUT[0]), .CK (clk), .D (n_0));
DFF_X1 \DATA_reg[1]  (.Q (DATA_OUT[1]), .CK (clk), .D (n_1));
DFF_X1 \DATA_reg[2]  (.Q (DATA_OUT[2]), .CK (clk), .D (n_2));
DFF_X1 \DATA_reg[3]  (.Q (DATA_OUT[3]), .CK (clk), .D (n_3));
DFF_X1 \DATA_reg[4]  (.Q (DATA_OUT[4]), .CK (clk), .D (n_4));
DFF_X1 \DATA_reg[5]  (.Q (DATA_OUT[5]), .CK (clk), .D (n_5));
DFF_X1 \DATA_reg[6]  (.Q (DATA_OUT[6]), .CK (clk), .D (n_6));
DFF_X1 \DATA_reg[7]  (.Q (DATA_OUT[7]), .CK (clk), .D (n_7));
DFF_X1 \DATA_reg[8]  (.Q (DATA_OUT[8]), .CK (clk), .D (n_8));
DFF_X1 \DATA_reg[9]  (.Q (DATA_OUT[9]), .CK (clk), .D (n_9));
DFF_X1 \DATA_reg[10]  (.Q (DATA_OUT[10]), .CK (clk), .D (n_10));
DFF_X1 \DATA_reg[11]  (.Q (DATA_OUT[11]), .CK (clk), .D (n_11));
DFF_X1 \DATA_reg[12]  (.Q (DATA_OUT[12]), .CK (clk), .D (n_12));
DFF_X1 \DATA_reg[13]  (.Q (DATA_OUT[13]), .CK (clk), .D (n_13));
DFF_X1 \DATA_reg[14]  (.Q (DATA_OUT[14]), .CK (clk), .D (n_14));
DFF_X1 \DATA_reg[15]  (.Q (DATA_OUT[15]), .CK (clk), .D (n_15));
DFF_X1 \DATA_reg[16]  (.Q (DATA_OUT[16]), .CK (clk), .D (n_16));
DFF_X1 \DATA_reg[17]  (.Q (DATA_OUT[17]), .CK (clk), .D (n_17));
DFF_X1 \DATA_reg[18]  (.Q (DATA_OUT[18]), .CK (clk), .D (n_18));
DFF_X1 \DATA_reg[19]  (.Q (DATA_OUT[19]), .CK (clk), .D (n_19));
DFF_X1 \DATA_reg[20]  (.Q (DATA_OUT[20]), .CK (clk), .D (n_20));
DFF_X1 \DATA_reg[21]  (.Q (DATA_OUT[21]), .CK (clk), .D (n_21));
DFF_X1 \DATA_reg[22]  (.Q (DATA_OUT[22]), .CK (clk), .D (n_22));
DFF_X1 \DATA_reg[23]  (.Q (DATA_OUT[23]), .CK (clk), .D (n_23));
DFF_X1 \DATA_reg[24]  (.Q (DATA_OUT[24]), .CK (clk), .D (n_24));
DFF_X1 \DATA_reg[25]  (.Q (DATA_OUT[25]), .CK (clk), .D (n_25));
DFF_X1 \DATA_reg[26]  (.Q (DATA_OUT[26]), .CK (clk), .D (n_26));
DFF_X1 \DATA_reg[27]  (.Q (DATA_OUT[27]), .CK (clk), .D (n_27));
DFF_X1 \DATA_reg[28]  (.Q (DATA_OUT[28]), .CK (clk), .D (n_28));
DFF_X1 \DATA_reg[29]  (.Q (DATA_OUT[29]), .CK (clk), .D (n_29));
DFF_X1 \DATA_reg[30]  (.Q (DATA_OUT[30]), .CK (clk), .D (n_30));
DFF_X1 \DATA_reg[31]  (.Q (DATA_OUT[31]), .CK (clk), .D (n_31));
DFF_X1 \DATA_reg[32]  (.Q (DATA_OUT[32]), .CK (clk), .D (n_32));
DFF_X1 \DATA_reg[33]  (.Q (DATA_OUT[33]), .CK (clk), .D (n_33));
DFF_X1 \DATA_reg[34]  (.Q (DATA_OUT[34]), .CK (clk), .D (n_34));
DFF_X1 \DATA_reg[35]  (.Q (DATA_OUT[35]), .CK (clk), .D (n_35));
DFF_X1 \DATA_reg[36]  (.Q (DATA_OUT[36]), .CK (clk), .D (n_36));
DFF_X1 \DATA_reg[37]  (.Q (DATA_OUT[37]), .CK (clk), .D (n_37));
DFF_X1 \DATA_reg[38]  (.Q (DATA_OUT[38]), .CK (clk), .D (n_38));
DFF_X1 \DATA_reg[39]  (.Q (DATA_OUT[39]), .CK (clk), .D (n_39));
DFF_X1 \DATA_reg[40]  (.Q (DATA_OUT[40]), .CK (clk), .D (n_40));
DFF_X1 \DATA_reg[41]  (.Q (DATA_OUT[41]), .CK (clk), .D (n_41));
DFF_X1 \DATA_reg[42]  (.Q (DATA_OUT[42]), .CK (clk), .D (n_42));
DFF_X1 \DATA_reg[43]  (.Q (DATA_OUT[43]), .CK (clk), .D (n_43));
DFF_X1 \DATA_reg[44]  (.Q (DATA_OUT[44]), .CK (clk), .D (n_44));
DFF_X1 \DATA_reg[45]  (.Q (DATA_OUT[45]), .CK (clk), .D (n_45));
DFF_X1 \DATA_reg[46]  (.Q (DATA_OUT[46]), .CK (clk), .D (n_46));
DFF_X1 \DATA_reg[47]  (.Q (DATA_OUT[47]), .CK (clk), .D (n_47));
DFF_X1 \DATA_reg[48]  (.Q (DATA_OUT[48]), .CK (clk), .D (n_48));
DFF_X1 \DATA_reg[49]  (.Q (DATA_OUT[49]), .CK (clk), .D (n_49));
DFF_X1 \DATA_reg[50]  (.Q (DATA_OUT[50]), .CK (clk), .D (n_50));
DFF_X1 \DATA_reg[51]  (.Q (DATA_OUT[51]), .CK (clk), .D (n_51));
DFF_X1 \DATA_reg[52]  (.Q (DATA_OUT[52]), .CK (clk), .D (n_52));
DFF_X1 \DATA_reg[53]  (.Q (DATA_OUT[53]), .CK (clk), .D (n_53));
DFF_X1 \DATA_reg[54]  (.Q (DATA_OUT[54]), .CK (clk), .D (n_54));
DFF_X1 \DATA_reg[55]  (.Q (DATA_OUT[55]), .CK (clk), .D (n_55));
DFF_X1 \DATA_reg[56]  (.Q (DATA_OUT[56]), .CK (clk), .D (n_56));
DFF_X1 \DATA_reg[57]  (.Q (DATA_OUT[57]), .CK (clk), .D (n_57));
DFF_X1 \DATA_reg[58]  (.Q (DATA_OUT[58]), .CK (clk), .D (n_58));
DFF_X1 \DATA_reg[59]  (.Q (DATA_OUT[59]), .CK (clk), .D (n_59));
DFF_X1 \DATA_reg[60]  (.Q (DATA_OUT[60]), .CK (clk), .D (n_60));
DFF_X1 \DATA_reg[61]  (.Q (DATA_OUT[61]), .CK (clk), .D (n_61));
DFF_X1 \DATA_reg[62]  (.Q (DATA_OUT[62]), .CK (clk), .D (n_62));
DFF_X1 \DATA_reg[63]  (.Q (DATA_OUT[63]), .CK (clk), .D (n_63));

endmodule //register__parameterized0

module register (DATA_IN, DATA_OUT, clk, reset);

output [31:0] DATA_OUT;
input [31:0] DATA_IN;
input clk;
input reset;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;
wire sps__n1;
wire spt__n3;


AND2_X1 i_0_31 (.ZN (n_31), .A1 (reset), .A2 (DATA_IN[31]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (reset), .A2 (DATA_IN[30]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (reset), .A2 (DATA_IN[29]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (reset), .A2 (DATA_IN[28]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (reset), .A2 (DATA_IN[27]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (reset), .A2 (DATA_IN[26]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (reset), .A2 (DATA_IN[25]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (reset), .A2 (DATA_IN[24]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (reset), .A2 (DATA_IN[23]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (reset), .A2 (DATA_IN[22]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (reset), .A2 (DATA_IN[21]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (reset), .A2 (DATA_IN[20]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (reset), .A2 (DATA_IN[19]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (reset), .A2 (DATA_IN[18]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (reset), .A2 (DATA_IN[17]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (reset), .A2 (DATA_IN[16]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (reset), .A2 (DATA_IN[15]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (reset), .A2 (DATA_IN[14]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (reset), .A2 (DATA_IN[13]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (reset), .A2 (DATA_IN[12]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (reset), .A2 (DATA_IN[11]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (reset), .A2 (DATA_IN[10]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (reset), .A2 (DATA_IN[9]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (reset), .A2 (DATA_IN[8]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (reset), .A2 (DATA_IN[7]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (reset), .A2 (DATA_IN[6]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (reset), .A2 (DATA_IN[5]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (reset), .A2 (DATA_IN[4]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (reset), .A2 (DATA_IN[3]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (reset), .A2 (DATA_IN[2]));
AND2_X1 i_0_1 (.ZN (n_1), .A1 (reset), .A2 (DATA_IN[1]));
AND2_X1 i_0_0 (.ZN (n_0), .A1 (DATA_IN[0]), .A2 (reset));
DFF_X1 \DATA_reg[0]  (.Q (spt__n3), .CK (clk), .D (n_0));
DFF_X1 \DATA_reg[1]  (.Q (DATA_OUT[1]), .CK (clk), .D (n_1));
DFF_X1 \DATA_reg[2]  (.Q (DATA_OUT[2]), .CK (clk), .D (n_2));
DFF_X1 \DATA_reg[3]  (.Q (DATA_OUT[3]), .CK (clk), .D (n_3));
DFF_X1 \DATA_reg[4]  (.Q (DATA_OUT[4]), .CK (clk), .D (n_4));
DFF_X1 \DATA_reg[5]  (.Q (DATA_OUT[5]), .CK (clk), .D (n_5));
DFF_X1 \DATA_reg[6]  (.Q (DATA_OUT[6]), .CK (clk), .D (n_6));
DFF_X1 \DATA_reg[7]  (.Q (DATA_OUT[7]), .CK (clk), .D (n_7));
DFF_X1 \DATA_reg[8]  (.Q (DATA_OUT[8]), .CK (clk), .D (n_8));
DFF_X1 \DATA_reg[9]  (.Q (DATA_OUT[9]), .CK (clk), .D (n_9));
DFF_X1 \DATA_reg[10]  (.Q (DATA_OUT[10]), .CK (clk), .D (n_10));
DFF_X1 \DATA_reg[11]  (.Q (DATA_OUT[11]), .CK (clk), .D (n_11));
DFF_X1 \DATA_reg[12]  (.Q (DATA_OUT[12]), .CK (clk), .D (n_12));
DFF_X1 \DATA_reg[13]  (.Q (DATA_OUT[13]), .CK (clk), .D (n_13));
DFF_X1 \DATA_reg[14]  (.Q (DATA_OUT[14]), .CK (clk), .D (n_14));
DFF_X1 \DATA_reg[15]  (.Q (DATA_OUT[15]), .CK (clk), .D (n_15));
DFF_X1 \DATA_reg[16]  (.Q (DATA_OUT[16]), .CK (clk), .D (n_16));
DFF_X1 \DATA_reg[17]  (.Q (DATA_OUT[17]), .CK (clk), .D (n_17));
DFF_X1 \DATA_reg[18]  (.Q (DATA_OUT[18]), .CK (clk), .D (n_18));
DFF_X1 \DATA_reg[19]  (.Q (DATA_OUT[19]), .CK (clk), .D (n_19));
DFF_X1 \DATA_reg[20]  (.Q (DATA_OUT[20]), .CK (clk), .D (n_20));
DFF_X1 \DATA_reg[21]  (.Q (DATA_OUT[21]), .CK (clk), .D (n_21));
DFF_X1 \DATA_reg[22]  (.Q (DATA_OUT[22]), .CK (clk), .D (n_22));
DFF_X1 \DATA_reg[23]  (.Q (DATA_OUT[23]), .CK (clk), .D (n_23));
DFF_X1 \DATA_reg[24]  (.Q (DATA_OUT[24]), .CK (clk), .D (n_24));
DFF_X1 \DATA_reg[25]  (.Q (DATA_OUT[25]), .CK (clk), .D (n_25));
DFF_X1 \DATA_reg[26]  (.Q (DATA_OUT[26]), .CK (clk), .D (n_26));
DFF_X1 \DATA_reg[27]  (.Q (DATA_OUT[27]), .CK (clk), .D (n_27));
DFF_X1 \DATA_reg[28]  (.Q (DATA_OUT[28]), .CK (clk), .D (n_28));
DFF_X1 \DATA_reg[29]  (.Q (DATA_OUT[29]), .CK (clk), .D (n_29));
DFF_X1 \DATA_reg[30]  (.Q (DATA_OUT[30]), .CK (clk), .D (n_30));
DFF_X1 \DATA_reg[31]  (.Q (sps__n1), .CK (clk), .D (n_31));
BUF_X8 sps__L1_c1_c1 (.Z (DATA_OUT[31]), .A (sps__n1));
BUF_X4 spt__c3 (.Z (DATA_OUT[0]), .A (spt__n3));

endmodule //register

module register__3_1 (DATA_IN, DATA_OUT, clk, reset);

output [31:0] DATA_OUT;
input [31:0] DATA_IN;
input clk;
input reset;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;
wire sps__n1;
wire spt__n3;


AND2_X1 i_0_31 (.ZN (n_31), .A1 (reset), .A2 (DATA_IN[31]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (reset), .A2 (DATA_IN[30]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (reset), .A2 (DATA_IN[29]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (reset), .A2 (DATA_IN[28]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (reset), .A2 (DATA_IN[27]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (reset), .A2 (DATA_IN[26]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (reset), .A2 (DATA_IN[25]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (reset), .A2 (DATA_IN[24]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (reset), .A2 (DATA_IN[23]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (reset), .A2 (DATA_IN[22]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (reset), .A2 (DATA_IN[21]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (reset), .A2 (DATA_IN[20]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (reset), .A2 (DATA_IN[19]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (reset), .A2 (DATA_IN[18]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (reset), .A2 (DATA_IN[17]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (reset), .A2 (DATA_IN[16]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (reset), .A2 (DATA_IN[15]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (reset), .A2 (DATA_IN[14]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (reset), .A2 (DATA_IN[13]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (reset), .A2 (DATA_IN[12]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (reset), .A2 (DATA_IN[11]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (reset), .A2 (DATA_IN[10]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (reset), .A2 (DATA_IN[9]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (reset), .A2 (DATA_IN[8]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (reset), .A2 (DATA_IN[7]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (reset), .A2 (DATA_IN[6]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (reset), .A2 (DATA_IN[5]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (reset), .A2 (DATA_IN[4]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (reset), .A2 (DATA_IN[3]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (reset), .A2 (DATA_IN[2]));
AND2_X1 i_0_1 (.ZN (n_1), .A1 (reset), .A2 (DATA_IN[1]));
AND2_X1 i_0_0 (.ZN (n_0), .A1 (DATA_IN[0]), .A2 (reset));
DFF_X1 \DATA_reg[0]  (.Q (spt__n3), .CK (clk), .D (n_0));
DFF_X1 \DATA_reg[1]  (.Q (DATA_OUT[1]), .CK (clk), .D (n_1));
DFF_X1 \DATA_reg[2]  (.Q (DATA_OUT[2]), .CK (clk), .D (n_2));
DFF_X1 \DATA_reg[3]  (.Q (DATA_OUT[3]), .CK (clk), .D (n_3));
DFF_X1 \DATA_reg[4]  (.Q (DATA_OUT[4]), .CK (clk), .D (n_4));
DFF_X1 \DATA_reg[5]  (.Q (DATA_OUT[5]), .CK (clk), .D (n_5));
DFF_X1 \DATA_reg[6]  (.Q (DATA_OUT[6]), .CK (clk), .D (n_6));
DFF_X1 \DATA_reg[7]  (.Q (DATA_OUT[7]), .CK (clk), .D (n_7));
DFF_X1 \DATA_reg[8]  (.Q (DATA_OUT[8]), .CK (clk), .D (n_8));
DFF_X1 \DATA_reg[9]  (.Q (DATA_OUT[9]), .CK (clk), .D (n_9));
DFF_X1 \DATA_reg[10]  (.Q (DATA_OUT[10]), .CK (clk), .D (n_10));
DFF_X1 \DATA_reg[11]  (.Q (DATA_OUT[11]), .CK (clk), .D (n_11));
DFF_X1 \DATA_reg[12]  (.Q (DATA_OUT[12]), .CK (clk), .D (n_12));
DFF_X1 \DATA_reg[13]  (.Q (DATA_OUT[13]), .CK (clk), .D (n_13));
DFF_X1 \DATA_reg[14]  (.Q (DATA_OUT[14]), .CK (clk), .D (n_14));
DFF_X1 \DATA_reg[15]  (.Q (DATA_OUT[15]), .CK (clk), .D (n_15));
DFF_X1 \DATA_reg[16]  (.Q (DATA_OUT[16]), .CK (clk), .D (n_16));
DFF_X1 \DATA_reg[17]  (.Q (DATA_OUT[17]), .CK (clk), .D (n_17));
DFF_X1 \DATA_reg[18]  (.Q (DATA_OUT[18]), .CK (clk), .D (n_18));
DFF_X1 \DATA_reg[19]  (.Q (DATA_OUT[19]), .CK (clk), .D (n_19));
DFF_X1 \DATA_reg[20]  (.Q (DATA_OUT[20]), .CK (clk), .D (n_20));
DFF_X1 \DATA_reg[21]  (.Q (DATA_OUT[21]), .CK (clk), .D (n_21));
DFF_X1 \DATA_reg[22]  (.Q (DATA_OUT[22]), .CK (clk), .D (n_22));
DFF_X1 \DATA_reg[23]  (.Q (DATA_OUT[23]), .CK (clk), .D (n_23));
DFF_X1 \DATA_reg[24]  (.Q (DATA_OUT[24]), .CK (clk), .D (n_24));
DFF_X1 \DATA_reg[25]  (.Q (DATA_OUT[25]), .CK (clk), .D (n_25));
DFF_X1 \DATA_reg[26]  (.Q (DATA_OUT[26]), .CK (clk), .D (n_26));
DFF_X1 \DATA_reg[27]  (.Q (DATA_OUT[27]), .CK (clk), .D (n_27));
DFF_X1 \DATA_reg[28]  (.Q (DATA_OUT[28]), .CK (clk), .D (n_28));
DFF_X1 \DATA_reg[29]  (.Q (DATA_OUT[29]), .CK (clk), .D (n_29));
DFF_X1 \DATA_reg[30]  (.Q (DATA_OUT[30]), .CK (clk), .D (n_30));
DFF_X1 \DATA_reg[31]  (.Q (sps__n1), .CK (clk), .D (n_31));
BUF_X8 sps__L1_c1_c1 (.Z (DATA_OUT[31]), .A (sps__n1));
BUF_X4 spt__c3 (.Z (DATA_OUT[0]), .A (spt__n3));

endmodule //register__3_1

module FA__2_140 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_140

module HA__2_374 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_374

module FA__2_137 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_137

module FA__2_134 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_134

module HA__2_371 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_371

module FA__2_131 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_131

module FA__2_128 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_128

module HA__2_368 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_368

module FA__2_125 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_125

module FA__2_122 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_122

module FA__2_119 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_119

module HA__2_365 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_365

module FA__2_116 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_116

module HA__2_362 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_362

module FA__2_113 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_113

module FA__2_110 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_110

module FA__2_107 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_107

module FA__2_104 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_104

module FA__2_101 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_101

module FA__2_98 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_98

module FA__2_95 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_95

module FA__2_92 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_92

module FA__2_89 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_89

module FA__2_86 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_86

module FA__2_83 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_83

module FA__2_80 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_80

module FA__2_77 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_77

module FA__2_74 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_74

module FA__2_71 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_71

module FA__2_68 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_68

module FA__2_65 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_65

module HA__2_359 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_359

module FA__2_62 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_62

module FA__2_59 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_59

module FA__2_56 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_56

module FA__2_53 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_53

module FA__2_50 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_50

module FA__2_47 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_47

module FA__2_44 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_44

module FA__2_41 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_41

module HA__2_356 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_356

module FA__2_38 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_38

module HA__2_353 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_353

module FA__2_35 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_35

module FA__2_32 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_32

module FA__2_29 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_29

module HA__2_350 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_350

module HA__2_347 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_347

module HA__2_344 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_344

module HA__2_341 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_341

module HA__2_338 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_338

module HA__2_335 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_335

module HA__2_332 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_332

module FA__2_26 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_26

module FA__2_23 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_23

module FA__2_20 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_20

module FA__2_17 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_17

module HA__2_329 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_329

module FA__2_14 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_14

module FA__2_11 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_11

module FA__2_8 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_8

module FA__2_5 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_5

module FA__2_2 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2

module WTM8 (A_7_PP_0, A_5_PP_0, B_7_PP_0, B_7_PP_1, B_7_PP_2, B_5_PP_0, B_5_PP_1, 
    B_5_PP_2, B_5_PP_3, A_7_PP_0PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_7_PP_0;
input A_5_PP_0;
input B_7_PP_0;
input B_7_PP_1;
input B_7_PP_2;
input B_5_PP_0;
input B_5_PP_1;
input B_5_PP_2;
input B_5_PP_3;
input A_7_PP_0PP_0;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A_7_PP_0PP_0), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A_5_PP_0), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A_7_PP_0PP_0), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A_5_PP_0), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A_7_PP_0), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A_5_PP_0), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A_5_PP_0), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A_5_PP_0), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A_5_PP_0), .A2 (B_5_PP_0));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B_5_PP_2));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B_5_PP_1));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B_5_PP_2));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B_5_PP_3));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B_5_PP_3));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B_7_PP_0));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B_7_PP_0));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B_7_PP_0));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B_7_PP_1));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B_7_PP_1));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B_7_PP_2));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_140 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_374 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_137 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_134 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_371 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_131 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_128 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_368 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_125 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_122 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_119 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_365 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_116 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_362 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_113 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_110 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_107 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_104 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_101 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_98 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_95 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_92 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_89 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_86 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_83 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_80 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_77 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_74 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_71 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_68 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_65 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_359 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_62 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_59 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_56 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_53 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_50 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_47 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_44 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_41 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_356 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_38 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_353 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_35 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_32 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_29 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_350 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_347 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_344 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_341 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_338 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_335 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_332 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_26 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_23 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_20 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_17 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_329 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_14 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_11 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_8 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_5 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_2 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8

module FA__2_1711 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_1711

module HA__2_1714 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1714

module FA__2_1717 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1717

module FA__2_1720 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1720

module HA__2_1723 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1723

module FA__2_1726 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1726

module FA__2_1729 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1729

module HA__2_1732 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1732

module FA__2_1735 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1735

module FA__2_1738 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1738

module FA__2_1741 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1741

module HA__2_1744 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1744

module FA__2_1747 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1747

module HA__2_1750 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1750

module FA__2_1753 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1753

module FA__2_1756 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1756

module FA__2_1759 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1759

module FA__2_1762 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1762

module FA__2_1765 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1765

module FA__2_1768 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1768

module FA__2_1771 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1771

module FA__2_1774 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1774

module FA__2_1777 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1777

module FA__2_1780 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1780

module FA__2_1783 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1783

module FA__2_1786 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1786

module FA__2_1789 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1789

module FA__2_1792 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1792

module FA__2_1795 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1795

module FA__2_1798 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1798

module FA__2_1801 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1801

module HA__2_1804 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1804

module FA__2_1807 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1807

module FA__2_1810 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1810

module FA__2_1813 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1813

module FA__2_1816 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1816

module FA__2_1819 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1819

module FA__2_1822 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1822

module FA__2_1825 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1825

module FA__2_1828 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1828

module HA__2_1831 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1831

module FA__2_1834 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1834

module HA__2_1837 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1837

module FA__2_1840 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1840

module FA__2_1843 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1843

module FA__2_1846 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1846

module HA__2_1849 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1849

module HA__2_1852 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1852

module HA__2_1855 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1855

module HA__2_1858 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1858

module HA__2_1861 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1861

module HA__2_1864 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1864

module HA__2_1867 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1867

module FA__2_1870 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1870

module FA__2_1873 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1873

module FA__2_1876 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1876

module FA__2_1879 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1879

module HA__2_1882 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1882

module FA__2_1885 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1885

module FA__2_1888 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1888

module FA__2_1891 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1891

module FA__2_1894 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1894

module FA__2_1897 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1897

module WTM8__2_1898 (A_5_PP_0, A_5_PP_1, A_4_PP_0, A_4_PP_1, A_4_PP_2, A_4_PP_3, 
    A_4_PP_4, B_5_PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_5_PP_0;
input A_5_PP_1;
input A_4_PP_0;
input A_4_PP_1;
input A_4_PP_2;
input A_4_PP_3;
input A_4_PP_4;
input B_5_PP_0;
wire spw_n83;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A_4_PP_3), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X4 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A_5_PP_1), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A_5_PP_1), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A_4_PP_4), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A_5_PP_0), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A_4_PP_2), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A_4_PP_1), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (spw_n83), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B_5_PP_0));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (spw_n83), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_1711 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_1714 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_1717 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_1720 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_1723 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_1726 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_1729 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_1732 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_1735 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_1738 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_1741 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_1744 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_1747 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_1750 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_1753 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_1756 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_1759 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_1762 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_1765 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_1768 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_1771 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_1774 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_1777 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_1780 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_1783 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_1786 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_1789 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_1792 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_1795 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_1798 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_1801 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_1804 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_1807 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_1810 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_1813 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_1816 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_1819 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_1822 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_1825 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_1828 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_1831 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_1834 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_1837 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_1840 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_1843 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_1846 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_1849 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_1852 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_1855 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_1858 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_1861 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_1864 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_1867 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_1870 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_1873 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_1876 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_1879 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_1882 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_1885 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_1888 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_1891 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_1894 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_1897 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));
BUF_X1 spw__L1_c3_c1 (.Z (spw_n83), .A (A_4_PP_0));

endmodule //WTM8__2_1898

module FA__2_1457 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_1457

module HA__2_1460 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1460

module FA__2_1463 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1463

module FA__2_1466 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1466

module HA__2_1469 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1469

module FA__2_1472 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1472

module FA__2_1475 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1475

module HA__2_1478 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1478

module FA__2_1481 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1481

module FA__2_1484 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1484

module FA__2_1487 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1487

module HA__2_1490 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1490

module FA__2_1493 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1493

module HA__2_1496 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1496

module FA__2_1499 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1499

module FA__2_1502 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1502

module FA__2_1505 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1505

module FA__2_1508 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1508

module FA__2_1511 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1511

module FA__2_1514 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1514

module FA__2_1517 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1517

module FA__2_1520 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1520

module FA__2_1523 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1523

module FA__2_1526 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1526

module FA__2_1529 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1529

module FA__2_1532 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1532

module FA__2_1535 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1535

module FA__2_1538 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1538

module FA__2_1541 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1541

module FA__2_1544 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1544

module FA__2_1547 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1547

module HA__2_1550 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1550

module FA__2_1553 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1553

module FA__2_1556 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1556

module FA__2_1559 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1559

module FA__2_1562 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1562

module FA__2_1565 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1565

module FA__2_1568 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1568

module FA__2_1571 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1571

module FA__2_1574 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1574

module HA__2_1577 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1577

module FA__2_1580 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1580

module HA__2_1583 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1583

module FA__2_1586 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1586

module FA__2_1589 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1589

module FA__2_1592 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1592

module HA__2_1595 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1595

module HA__2_1598 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1598

module HA__2_1601 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1601

module HA__2_1604 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1604

module HA__2_1607 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1607

module HA__2_1610 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1610

module HA__2_1613 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1613

module FA__2_1616 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1616

module FA__2_1619 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1619

module FA__2_1622 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1622

module FA__2_1625 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1625

module HA__2_1628 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1628

module FA__2_1631 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1631

module FA__2_1634 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1634

module FA__2_1637 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1637

module FA__2_1640 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1640

module FA__2_1643 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1643

module WTM8__2_1644 (A_4_PP_0, B_7_PP_0, B_7_PP_1, A_6_PP_0, A_6_PP_1, A_6_PP_2, 
    A_6_PP_3, A_7_PP_0, A_7_PP_1, B_5_PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_4_PP_0;
input B_7_PP_0;
input B_7_PP_1;
input A_6_PP_0;
input A_6_PP_1;
input A_6_PP_2;
input A_6_PP_3;
input A_7_PP_0;
input A_7_PP_1;
input B_5_PP_0;
wire spw_n30;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;
wire spw__n12;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A_6_PP_0), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (spw_n30), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A_7_PP_0), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A_6_PP_3), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A_6_PP_2), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A_7_PP_1), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A_6_PP_1), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A_6_PP_1), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (spw__n12), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A_6_PP_1), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (spw_n30), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A_6_PP_0), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B_5_PP_0));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (spw_n30), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B_5_PP_0));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B_5_PP_0));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B_5_PP_0));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B_7_PP_0));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B_7_PP_0));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (spw_n30), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B_7_PP_0));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B_7_PP_0));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B_7_PP_1));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_1457 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_1460 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_1463 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_1466 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_1469 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_1472 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_1475 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_1478 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_1481 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_1484 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_1487 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_1490 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_1493 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_1496 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_1499 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_1502 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_1505 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_1508 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_1511 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_1514 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_1517 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_1520 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_1523 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_1526 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_1529 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_1532 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_1535 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_1538 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_1541 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_1544 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_1547 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_1550 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_1553 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_1556 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_1559 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_1562 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_1565 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_1568 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_1571 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_1574 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_1577 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_1580 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_1583 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_1586 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_1589 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_1592 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_1595 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_1598 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_1601 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_1604 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_1607 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_1610 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_1613 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_1616 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_1619 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_1622 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_1625 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_1628 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_1631 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_1634 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_1637 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_1640 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_1643 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));
BUF_X2 spw__L3_c6_c1 (.Z (spw_n30), .A (spw__n12));
BUF_X1 spw__L2_c5_c2 (.Z (spw__n12), .A (A_4_PP_0));

endmodule //WTM8__2_1644

module FA__2_257 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_257

module FA__2_254 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_254

module FA__2_251 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_251

module FA__2_248 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_248

module FA__2_245 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_245

module FA__2_242 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_242

module FA__2_239 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X2 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_239

module FA__2_236 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_236

module FA__2_233 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_233

module FA__2_230 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_230

module FA__2_227 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_227

module FA__2_224 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_224

module FA__2_221 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_221

module FA__2_218 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_218

module FA__2_215 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_215

module FA__2_212 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_212

module adder64 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;


FA__2_257 genblk1_39_F (.carry (z[40]), .sum (z[39]), .b (y[39]), .cin (\carry[38] ));
FA__2_254 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .b (y[38]), .cin (\carry[37] ));
FA__2_251 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .b (y[37]), .cin (\carry[36] ));
FA__2_248 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .b (y[36]), .cin (\carry[35] ));
FA__2_245 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .b (y[35]), .cin (\carry[34] ));
FA__2_242 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .b (y[34]), .cin (\carry[33] ));
FA__2_239 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .b (y[33]), .cin (\carry[32] ));
FA__2_236 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .b (y[32]), .cin (\carry[31] ));
FA__2_233 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .a (x[31]), .b (y[31]), .cin (\carry[30] ));
FA__2_230 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .a (x[30]), .b (y[30]), .cin (\carry[29] ));
FA__2_227 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .a (x[29]), .b (y[29])
    , .cin (\carry[28] ));
FA__2_224 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .a (x[28]), .b (y[28]), .cin (\carry[27] ));
FA__2_221 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .a (x[27]), .b (y[27]), .cin (\carry[26] ));
FA__2_218 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .a (x[26]), .b (y[26]), .cin (\carry[25] ));
FA__2_215 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .a (x[25]), .b (y[25])
    , .cin (\carry[24] ));
FA__2_212 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24]));

endmodule //adder64

module FA__2_1203 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_1203

module HA__2_1206 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1206

module FA__2_1209 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1209

module FA__2_1212 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1212

module HA__2_1215 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1215

module FA__2_1218 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1218

module FA__2_1221 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1221

module HA__2_1224 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1224

module FA__2_1227 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1227

module FA__2_1230 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1230

module FA__2_1233 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1233

module HA__2_1236 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1236

module FA__2_1239 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1239

module HA__2_1242 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1242

module FA__2_1245 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1245

module FA__2_1248 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1248

module FA__2_1251 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1251

module FA__2_1254 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1254

module FA__2_1257 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1257

module FA__2_1260 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1260

module FA__2_1263 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1263

module FA__2_1266 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1266

module FA__2_1269 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1269

module FA__2_1272 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1272

module FA__2_1275 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1275

module FA__2_1278 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1278

module FA__2_1281 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1281

module FA__2_1284 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1284

module FA__2_1287 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1287

module FA__2_1290 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1290

module FA__2_1293 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1293

module HA__2_1296 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1296

module FA__2_1299 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1299

module FA__2_1302 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1302

module FA__2_1305 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1305

module FA__2_1308 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1308

module FA__2_1311 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1311

module FA__2_1314 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1314

module FA__2_1317 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1317

module FA__2_1320 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1320

module HA__2_1323 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1323

module FA__2_1326 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1326

module HA__2_1329 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1329

module FA__2_1332 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1332

module FA__2_1335 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1335

module FA__2_1338 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1338

module HA__2_1341 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1341

module HA__2_1344 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1344

module HA__2_1347 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1347

module HA__2_1350 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1350

module HA__2_1353 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1353

module HA__2_1356 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1356

module HA__2_1359 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1359

module FA__2_1362 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1362

module FA__2_1365 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1365

module FA__2_1368 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1368

module FA__2_1371 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1371

module HA__2_1374 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1374

module FA__2_1377 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1377

module FA__2_1380 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1380

module FA__2_1383 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1383

module FA__2_1386 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1386

module FA__2_1389 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1389

module WTM8__2_1390 (A_4_PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_4_PP_0;
wire spw_n8;
wire spw_n16;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (spw_n8), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (spw_n16), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A_4_PP_0), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (spw_n16), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (spw_n16), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A_4_PP_0), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (spw_n16), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (spw_n16), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (spw_n8), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (spw_n16), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (spw_n8), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (spw_n16), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (spw_n8), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (spw_n16), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_1203 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_1206 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_1209 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_1212 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_1215 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_1218 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_1221 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_1224 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_1227 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_1230 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_1233 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_1236 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_1239 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_1242 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_1245 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_1248 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_1251 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_1254 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_1257 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_1260 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_1263 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_1266 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_1269 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_1272 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_1275 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_1278 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_1281 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_1284 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_1287 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_1290 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_1293 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_1296 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_1299 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_1302 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_1305 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_1308 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_1311 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_1314 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_1317 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_1320 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_1323 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_1326 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_1329 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_1332 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_1335 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_1338 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_1341 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_1344 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_1347 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_1350 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_1353 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_1356 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_1359 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_1362 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_1365 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_1368 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_1371 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_1374 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_1377 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_1380 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_1383 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_1386 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_1389 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));
BUF_X1 spw__L4_c4_c1 (.Z (spw_n8), .A (A[5]));
BUF_X2 spw__L4_c4_c4 (.Z (spw_n16), .A (A[3]));

endmodule //WTM8__2_1390

module FA__2_2890 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2890

module FA__2_2893 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2893

module FA__2_2896 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2896

module FA__2_2899 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2899

module FA__2_2902 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2902

module FA__2_2905 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2905

module FA__2_2908 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2908

module FA__2_2911 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2911

module FA__2_2914 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2914

module FA__2_2917 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2917

module FA__2_2920 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2920

module FA__2_2923 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2923

module FA__2_2926 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2926

module FA__2_2929 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2929

module FA__2_2932 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2932

module FA__2_2935 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_2935

module adder64__2_3056 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;


FA__2_2890 genblk1_55_F (.carry (z[56]), .sum (z[55]), .b (y[55]), .cin (\carry[54] ));
FA__2_2893 genblk1_54_F (.carry (\carry[54] ), .sum (z[54]), .b (y[54]), .cin (\carry[53] ));
FA__2_2896 genblk1_53_F (.carry (\carry[53] ), .sum (z[53]), .b (y[53]), .cin (\carry[52] ));
FA__2_2899 genblk1_52_F (.carry (\carry[52] ), .sum (z[52]), .b (y[52]), .cin (\carry[51] ));
FA__2_2902 genblk1_51_F (.carry (\carry[51] ), .sum (z[51]), .b (y[51]), .cin (\carry[50] ));
FA__2_2905 genblk1_50_F (.carry (\carry[50] ), .sum (z[50]), .b (y[50]), .cin (\carry[49] ));
FA__2_2908 genblk1_49_F (.carry (\carry[49] ), .sum (z[49]), .b (y[49]), .cin (\carry[48] ));
FA__2_2911 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .b (y[48]), .cin (\carry[47] ));
FA__2_2914 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .a (x[47]), .b (y[47]), .cin (\carry[46] ));
FA__2_2917 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .a (x[46]), .b (y[46]), .cin (\carry[45] ));
FA__2_2920 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .a (x[45]), .b (y[45]), .cin (\carry[44] ));
FA__2_2923 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .a (x[44]), .b (y[44]), .cin (\carry[43] ));
FA__2_2926 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .a (x[43]), .b (y[43]), .cin (\carry[42] ));
FA__2_2929 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .a (x[42]), .b (y[42]), .cin (\carry[41] ));
FA__2_2932 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .a (x[41]), .b (y[41]), .cin (\carry[40] ));
FA__2_2935 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .a (x[40]), .b (y[40]));

endmodule //adder64__2_3056

module FA__2_2694 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2694

module FA__2_2697 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2697

module FA__2_2700 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2700

module FA__2_2703 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2703

module FA__2_2706 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2706

module FA__2_2709 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2709

module FA__2_2712 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2712

module FA__2_2715 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2715

module FA__2_2718 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2718

module FA__2_2721 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2721

module FA__2_2724 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2724

module FA__2_2727 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2727

module FA__2_2730 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2730

module FA__2_2733 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2733

module FA__2_2736 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2736

module FA__2_2739 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2739

module FA__2_2742 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2742

module FA__2_2745 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2745

module FA__2_2748 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2748

module FA__2_2751 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2751

module FA__2_2754 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2754

module FA__2_2757 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2757

module FA__2_2760 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2760

module FA__2_2763 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2763

module FA__2_2766 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_2766

module adder64__2_2863 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[55] ;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;


FA__2_2694 genblk1_56_F (.carry (z[57]), .sum (z[56]), .b (y[56]), .cin (\carry[55] ));
FA__2_2697 genblk1_55_F (.carry (\carry[55] ), .sum (z[55]), .b (y[55]), .cin (\carry[54] ));
FA__2_2700 genblk1_54_F (.carry (\carry[54] ), .sum (z[54]), .b (y[54]), .cin (\carry[53] ));
FA__2_2703 genblk1_53_F (.carry (\carry[53] ), .sum (z[53]), .b (y[53]), .cin (\carry[52] ));
FA__2_2706 genblk1_52_F (.carry (\carry[52] ), .sum (z[52]), .b (y[52]), .cin (\carry[51] ));
FA__2_2709 genblk1_51_F (.carry (\carry[51] ), .sum (z[51]), .b (y[51]), .cin (\carry[50] ));
FA__2_2712 genblk1_50_F (.carry (\carry[50] ), .sum (z[50]), .b (y[50]), .cin (\carry[49] ));
FA__2_2715 genblk1_49_F (.carry (\carry[49] ), .sum (z[49]), .b (y[49]), .cin (\carry[48] ));
FA__2_2718 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .b (y[48]), .cin (\carry[47] ));
FA__2_2721 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .b (y[47]), .cin (\carry[46] ));
FA__2_2724 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .b (y[46]), .cin (\carry[45] ));
FA__2_2727 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .b (y[45]), .cin (\carry[44] ));
FA__2_2730 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .b (y[44]), .cin (\carry[43] ));
FA__2_2733 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .b (y[43]), .cin (\carry[42] ));
FA__2_2736 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .b (y[42]), .cin (\carry[41] ));
FA__2_2739 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .b (y[41]), .cin (\carry[40] ));
FA__2_2742 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .a (x[40]), .b (y[40]), .cin (\carry[39] ));
FA__2_2745 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .a (x[39]), .b (y[39]), .cin (\carry[38] ));
FA__2_2748 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .a (x[38]), .b (y[38]), .cin (\carry[37] ));
FA__2_2751 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .a (x[37]), .b (y[37]), .cin (\carry[36] ));
FA__2_2754 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .a (x[36]), .b (y[36]), .cin (\carry[35] ));
FA__2_2757 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .a (x[35]), .b (y[35]), .cin (\carry[34] ));
FA__2_2760 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .a (x[34]), .b (y[34]), .cin (\carry[33] ));
FA__2_2763 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .a (x[33]), .b (y[33])
    , .cin (\carry[32] ));
FA__2_2766 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32]));

endmodule //adder64__2_2863

module FA__2_949 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_949

module HA__2_952 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_952

module FA__2_955 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_955

module FA__2_958 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_958

module HA__2_961 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_961

module FA__2_964 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_964

module FA__2_967 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_967

module HA__2_970 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_970

module FA__2_973 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_973

module FA__2_976 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_976

module FA__2_979 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_979

module HA__2_982 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_982

module FA__2_985 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_985

module HA__2_988 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_988

module FA__2_991 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_991

module FA__2_994 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_994

module FA__2_997 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_997

module FA__2_1000 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1000

module FA__2_1003 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1003

module FA__2_1006 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1006

module FA__2_1009 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1009

module FA__2_1012 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1012

module FA__2_1015 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1015

module FA__2_1018 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1018

module FA__2_1021 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1021

module FA__2_1024 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1024

module FA__2_1027 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1027

module FA__2_1030 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1030

module FA__2_1033 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1033

module FA__2_1036 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1036

module FA__2_1039 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1039

module HA__2_1042 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1042

module FA__2_1045 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1045

module FA__2_1048 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1048

module FA__2_1051 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1051

module FA__2_1054 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1054

module FA__2_1057 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1057

module FA__2_1060 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1060

module FA__2_1063 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1063

module FA__2_1066 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1066

module HA__2_1069 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1069

module FA__2_1072 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1072

module HA__2_1075 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1075

module FA__2_1078 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1078

module FA__2_1081 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1081

module FA__2_1084 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1084

module HA__2_1087 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1087

module HA__2_1090 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1090

module HA__2_1093 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1093

module HA__2_1096 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1096

module HA__2_1099 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1099

module HA__2_1102 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1102

module HA__2_1105 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1105

module FA__2_1108 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1108

module FA__2_1111 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1111

module FA__2_1114 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1114

module FA__2_1117 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1117

module HA__2_1120 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_1120

module FA__2_1123 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1123

module FA__2_1126 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1126

module FA__2_1129 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1129

module FA__2_1132 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1132

module FA__2_1135 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1135

module WTM8__2_1136 (A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_949 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_952 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_955 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_958 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_961 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_964 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_967 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_970 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_973 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_976 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_979 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_982 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_985 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_988 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_991 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_994 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_997 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_1000 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_1003 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_1006 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_1009 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_1012 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_1015 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_1018 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_1021 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_1024 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_1027 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_1030 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_1033 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_1036 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_1039 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_1042 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_1045 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_1048 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_1051 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_1054 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_1057 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_1060 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_1063 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_1066 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_1069 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_1072 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_1075 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_1078 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_1081 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_1084 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_1087 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_1090 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_1093 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_1096 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_1099 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_1102 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_1105 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_1108 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_1111 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_1114 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_1117 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_1120 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_1123 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_1126 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_1129 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_1132 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_1135 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__2_1136

module FA__2_2480 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


XOR2_X1 i_0_0 (.Z (sum), .A (b), .B (cin));

endmodule //FA__2_2480

module FA__2_2483 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2483

module FA__2_2486 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2486

module FA__2_2489 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2489

module FA__2_2492 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2492

module FA__2_2495 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2495

module FA__2_2498 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2498

module FA__2_2501 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2501

module FA__2_2504 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2504

module FA__2_2507 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2507

module FA__2_2510 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2510

module FA__2_2513 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2513

module FA__2_2516 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2516

module FA__2_2519 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2519

module FA__2_2522 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2522

module FA__2_2525 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2525

module FA__2_2528 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2528

module FA__2_2531 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2531

module FA__2_2534 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2534

module FA__2_2537 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2537

module FA__2_2540 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2540

module FA__2_2543 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2543

module FA__2_2546 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2546

module FA__2_2549 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2549

module FA__2_2552 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2552

module FA__2_2555 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2555

module FA__2_2558 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2558

module FA__2_2561 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2561

module FA__2_2564 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2564

module FA__2_2567 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2567

module FA__2_2570 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2570

module FA__2_2573 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2573

module FA__2_2576 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2576

module FA__2_2579 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2579

module FA__2_2582 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2582

module FA__2_2585 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2585

module FA__2_2588 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2588

module FA__2_2591 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2591

module FA__2_2594 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2594

module FA__2_2597 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_2597

module adder64__2_2670 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[62] ;
wire \carry[61] ;
wire \carry[60] ;
wire \carry[59] ;
wire \carry[58] ;
wire \carry[57] ;
wire \carry[56] ;
wire \carry[55] ;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;


FA__2_2480 genblk1_63_F (.sum (z[63]), .b (y[63]), .cin (\carry[62] ));
FA__2_2483 genblk1_62_F (.carry (\carry[62] ), .sum (z[62]), .b (y[62]), .cin (\carry[61] ));
FA__2_2486 genblk1_61_F (.carry (\carry[61] ), .sum (z[61]), .b (y[61]), .cin (\carry[60] ));
FA__2_2489 genblk1_60_F (.carry (\carry[60] ), .sum (z[60]), .b (y[60]), .cin (\carry[59] ));
FA__2_2492 genblk1_59_F (.carry (\carry[59] ), .sum (z[59]), .b (y[59]), .cin (\carry[58] ));
FA__2_2495 genblk1_58_F (.carry (\carry[58] ), .sum (z[58]), .b (y[58]), .cin (\carry[57] ));
FA__2_2498 genblk1_57_F (.carry (\carry[57] ), .sum (z[57]), .a (x[57]), .b (y[57]), .cin (\carry[56] ));
FA__2_2501 genblk1_56_F (.carry (\carry[56] ), .sum (z[56]), .a (x[56]), .b (y[56]), .cin (\carry[55] ));
FA__2_2504 genblk1_55_F (.carry (\carry[55] ), .sum (z[55]), .a (x[55]), .b (y[55]), .cin (\carry[54] ));
FA__2_2507 genblk1_54_F (.carry (\carry[54] ), .sum (z[54]), .a (x[54]), .b (y[54]), .cin (\carry[53] ));
FA__2_2510 genblk1_53_F (.carry (\carry[53] ), .sum (z[53]), .a (x[53]), .b (y[53]), .cin (\carry[52] ));
FA__2_2513 genblk1_52_F (.carry (\carry[52] ), .sum (z[52]), .a (x[52]), .b (y[52]), .cin (\carry[51] ));
FA__2_2516 genblk1_51_F (.carry (\carry[51] ), .sum (z[51]), .a (x[51]), .b (y[51]), .cin (\carry[50] ));
FA__2_2519 genblk1_50_F (.carry (\carry[50] ), .sum (z[50]), .a (x[50]), .b (y[50]), .cin (\carry[49] ));
FA__2_2522 genblk1_49_F (.carry (\carry[49] ), .sum (z[49]), .a (x[49]), .b (y[49]), .cin (\carry[48] ));
FA__2_2525 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .a (x[48]), .b (y[48]), .cin (\carry[47] ));
FA__2_2528 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .a (x[47]), .b (y[47]), .cin (\carry[46] ));
FA__2_2531 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .a (x[46]), .b (y[46]), .cin (\carry[45] ));
FA__2_2534 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .a (x[45]), .b (y[45]), .cin (\carry[44] ));
FA__2_2537 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .a (x[44]), .b (y[44]), .cin (\carry[43] ));
FA__2_2540 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .a (x[43]), .b (y[43]), .cin (\carry[42] ));
FA__2_2543 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .a (x[42]), .b (y[42]), .cin (\carry[41] ));
FA__2_2546 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .a (x[41]), .b (y[41]), .cin (\carry[40] ));
FA__2_2549 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .a (x[40]), .b (y[40])
    , .cin (\carry[39] ));
FA__2_2552 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .a (x[39]), .b (y[39])
    , .cin (\carry[38] ));
FA__2_2555 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .a (x[38]), .b (y[38]), .cin (\carry[37] ));
FA__2_2558 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .a (x[37]), .b (y[37])
    , .cin (\carry[36] ));
FA__2_2561 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .a (x[36]), .b (y[36]), .cin (\carry[35] ));
FA__2_2564 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .a (x[35]), .b (y[35])
    , .cin (\carry[34] ));
FA__2_2567 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .a (x[34]), .b (y[34])
    , .cin (\carry[33] ));
FA__2_2570 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .a (x[33]), .b (y[33]), .cin (\carry[32] ));
FA__2_2573 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32]), .cin (\carry[31] ));
FA__2_2576 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .a (x[31]), .b (y[31]), .cin (\carry[30] ));
FA__2_2579 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .a (x[30]), .b (y[30]), .cin (\carry[29] ));
FA__2_2582 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .a (x[29]), .b (y[29]), .cin (\carry[28] ));
FA__2_2585 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .a (x[28]), .b (y[28]), .cin (\carry[27] ));
FA__2_2588 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .a (x[27]), .b (y[27]), .cin (\carry[26] ));
FA__2_2591 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .a (x[26]), .b (y[26]), .cin (\carry[25] ));
FA__2_2594 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .a (x[25]), .b (y[25]), .cin (\carry[24] ));
FA__2_2597 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24]));

endmodule //adder64__2_2670

module FA__2_2287 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


XOR2_X1 i_0_0 (.Z (sum), .A (b), .B (cin));

endmodule //FA__2_2287

module FA__2_2290 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2290

module FA__2_2293 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2293

module FA__2_2296 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2296

module FA__2_2299 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2299

module FA__2_2302 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2302

module FA__2_2305 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2305

module FA__2_2308 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2308

module FA__2_2311 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2311

module FA__2_2314 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2314

module FA__2_2317 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2317

module FA__2_2320 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2320

module FA__2_2323 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2323

module FA__2_2326 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2326

module FA__2_2329 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2329

module FA__2_2332 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2332

module FA__2_2335 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2335

module FA__2_2338 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2338

module FA__2_2341 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2341

module FA__2_2344 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2344

module FA__2_2347 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2347

module FA__2_2350 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2350

module FA__2_2353 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2353

module FA__2_2356 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_2356

module adder64__2_2477 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[62] ;
wire \carry[61] ;
wire \carry[60] ;
wire \carry[59] ;
wire \carry[58] ;
wire \carry[57] ;
wire \carry[56] ;
wire \carry[55] ;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;


FA__2_2287 genblk1_63_F (.sum (z[63]), .b (y[63]), .cin (\carry[62] ));
FA__2_2290 genblk1_62_F (.carry (\carry[62] ), .sum (z[62]), .b (y[62]), .cin (\carry[61] ));
FA__2_2293 genblk1_61_F (.carry (\carry[61] ), .sum (z[61]), .b (y[61]), .cin (\carry[60] ));
FA__2_2296 genblk1_60_F (.carry (\carry[60] ), .sum (z[60]), .b (y[60]), .cin (\carry[59] ));
FA__2_2299 genblk1_59_F (.carry (\carry[59] ), .sum (z[59]), .b (y[59]), .cin (\carry[58] ));
FA__2_2302 genblk1_58_F (.carry (\carry[58] ), .sum (z[58]), .b (y[58]), .cin (\carry[57] ));
FA__2_2305 genblk1_57_F (.carry (\carry[57] ), .sum (z[57]), .b (y[57]), .cin (\carry[56] ));
FA__2_2308 genblk1_56_F (.carry (\carry[56] ), .sum (z[56]), .b (y[56]), .cin (\carry[55] ));
FA__2_2311 genblk1_55_F (.carry (\carry[55] ), .sum (z[55]), .b (y[55]), .cin (\carry[54] ));
FA__2_2314 genblk1_54_F (.carry (\carry[54] ), .sum (z[54]), .b (y[54]), .cin (\carry[53] ));
FA__2_2317 genblk1_53_F (.carry (\carry[53] ), .sum (z[53]), .b (y[53]), .cin (\carry[52] ));
FA__2_2320 genblk1_52_F (.carry (\carry[52] ), .sum (z[52]), .b (y[52]), .cin (\carry[51] ));
FA__2_2323 genblk1_51_F (.carry (\carry[51] ), .sum (z[51]), .b (y[51]), .cin (\carry[50] ));
FA__2_2326 genblk1_50_F (.carry (\carry[50] ), .sum (z[50]), .b (y[50]), .cin (\carry[49] ));
FA__2_2329 genblk1_49_F (.carry (\carry[49] ), .sum (z[49]), .b (y[49]), .cin (\carry[48] ));
FA__2_2332 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .a (x[48]), .b (y[48]), .cin (\carry[47] ));
FA__2_2335 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .a (x[47]), .b (y[47]), .cin (\carry[46] ));
FA__2_2338 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .a (x[46]), .b (y[46]), .cin (\carry[45] ));
FA__2_2341 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .a (x[45]), .b (y[45]), .cin (\carry[44] ));
FA__2_2344 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .a (x[44]), .b (y[44]), .cin (\carry[43] ));
FA__2_2347 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .a (x[43]), .b (y[43]), .cin (\carry[42] ));
FA__2_2350 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .a (x[42]), .b (y[42]), .cin (\carry[41] ));
FA__2_2353 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .a (x[41]), .b (y[41]), .cin (\carry[40] ));
FA__2_2356 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .a (x[40]), .b (y[40]));

endmodule //adder64__2_2477

module FA__2_2094 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


XOR2_X1 i_0_0 (.Z (sum), .A (b), .B (cin));

endmodule //FA__2_2094

module FA__2_2097 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2097

module FA__2_2100 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2100

module FA__2_2103 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2103

module FA__2_2106 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2106

module FA__2_2109 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2109

module FA__2_2112 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2112

module FA__2_2115 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_2115

module FA__2_2118 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2118

module FA__2_2121 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2121

module FA__2_2124 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2124

module FA__2_2127 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2127

module FA__2_2130 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2130

module FA__2_2133 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2133

module FA__2_2136 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_2136

module FA__2_2139 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_2139

module adder64__2_2284 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[62] ;
wire \carry[61] ;
wire \carry[60] ;
wire \carry[59] ;
wire \carry[58] ;
wire \carry[57] ;
wire \carry[56] ;
wire \carry[55] ;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;


FA__2_2094 genblk1_63_F (.sum (z[63]), .b (y[63]), .cin (\carry[62] ));
FA__2_2097 genblk1_62_F (.carry (\carry[62] ), .sum (z[62]), .b (y[62]), .cin (\carry[61] ));
FA__2_2100 genblk1_61_F (.carry (\carry[61] ), .sum (z[61]), .b (y[61]), .cin (\carry[60] ));
FA__2_2103 genblk1_60_F (.carry (\carry[60] ), .sum (z[60]), .b (y[60]), .cin (\carry[59] ));
FA__2_2106 genblk1_59_F (.carry (\carry[59] ), .sum (z[59]), .b (y[59]), .cin (\carry[58] ));
FA__2_2109 genblk1_58_F (.carry (\carry[58] ), .sum (z[58]), .b (y[58]), .cin (\carry[57] ));
FA__2_2112 genblk1_57_F (.carry (\carry[57] ), .sum (z[57]), .b (y[57]), .cin (\carry[56] ));
FA__2_2115 genblk1_56_F (.carry (\carry[56] ), .sum (z[56]), .b (y[56]), .cin (\carry[55] ));
FA__2_2118 genblk1_55_F (.carry (\carry[55] ), .sum (z[55]), .a (x[55]), .b (y[55]), .cin (\carry[54] ));
FA__2_2121 genblk1_54_F (.carry (\carry[54] ), .sum (z[54]), .a (x[54]), .b (y[54]), .cin (\carry[53] ));
FA__2_2124 genblk1_53_F (.carry (\carry[53] ), .sum (z[53]), .a (x[53]), .b (y[53]), .cin (\carry[52] ));
FA__2_2127 genblk1_52_F (.carry (\carry[52] ), .sum (z[52]), .a (x[52]), .b (y[52]), .cin (\carry[51] ));
FA__2_2130 genblk1_51_F (.carry (\carry[51] ), .sum (z[51]), .a (x[51]), .b (y[51]), .cin (\carry[50] ));
FA__2_2133 genblk1_50_F (.carry (\carry[50] ), .sum (z[50]), .a (x[50]), .b (y[50]), .cin (\carry[49] ));
FA__2_2136 genblk1_49_F (.carry (\carry[49] ), .sum (z[49]), .a (x[49]), .b (y[49]), .cin (\carry[48] ));
FA__2_2139 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .a (x[48]), .b (y[48]));

endmodule //adder64__2_2284

module FA__2_695 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_695

module HA__2_698 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_698

module FA__2_701 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_701

module FA__2_704 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_704

module HA__2_707 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_707

module FA__2_710 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_710

module FA__2_713 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_713

module HA__2_716 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_716

module FA__2_719 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_719

module FA__2_722 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_722

module FA__2_725 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_725

module HA__2_728 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_728

module FA__2_731 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_731

module HA__2_734 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_734

module FA__2_737 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_737

module FA__2_740 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_740

module FA__2_743 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_743

module FA__2_746 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_746

module FA__2_749 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_749

module FA__2_752 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_752

module FA__2_755 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_755

module FA__2_758 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_758

module FA__2_761 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_761

module FA__2_764 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_764

module FA__2_767 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_767

module FA__2_770 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_770

module FA__2_773 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_773

module FA__2_776 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_776

module FA__2_779 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_779

module FA__2_782 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_782

module FA__2_785 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_785

module HA__2_788 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_788

module FA__2_791 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_791

module FA__2_794 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_794

module FA__2_797 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_797

module FA__2_800 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_800

module FA__2_803 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_803

module FA__2_806 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_806

module FA__2_809 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_809

module FA__2_812 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_812

module HA__2_815 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_815

module FA__2_818 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_818

module HA__2_821 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_821

module FA__2_824 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_824

module FA__2_827 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_827

module FA__2_830 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_830

module HA__2_833 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_833

module HA__2_836 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_836

module HA__2_839 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_839

module HA__2_842 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_842

module HA__2_845 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_845

module HA__2_848 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_848

module HA__2_851 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_851

module FA__2_854 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_854

module FA__2_857 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_857

module FA__2_860 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_860

module FA__2_863 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_863

module HA__2_866 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_866

module FA__2_869 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_869

module FA__2_872 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_872

module FA__2_875 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_875

module FA__2_878 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_878

module FA__2_881 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_881

module WTM8__2_882 (A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_695 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_698 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_701 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_704 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_707 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_710 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_713 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_716 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_719 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_722 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_725 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_728 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_731 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_734 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_737 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_740 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_743 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_746 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_749 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_752 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_755 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_758 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_761 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_764 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_767 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_770 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_773 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_776 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_779 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_782 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_785 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_788 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_791 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_794 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_797 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_800 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_803 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_806 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_809 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_812 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_815 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_818 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_821 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_824 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_827 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_830 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_833 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_836 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_839 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_842 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_845 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_848 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_851 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_854 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_857 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_860 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_863 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_866 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_869 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_872 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_875 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_878 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_881 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__2_882

module FA__2_441 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__2_441

module HA__2_444 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_444

module FA__2_447 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_447

module FA__2_450 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_450

module HA__2_453 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_453

module FA__2_456 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_456

module FA__2_459 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_459

module HA__2_462 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_462

module FA__2_465 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_465

module FA__2_468 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_468

module FA__2_471 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_471

module HA__2_474 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_474

module FA__2_477 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_477

module HA__2_480 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_480

module FA__2_483 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_483

module FA__2_486 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_486

module FA__2_489 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_489

module FA__2_492 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_492

module FA__2_495 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_495

module FA__2_498 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_498

module FA__2_501 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_501

module FA__2_504 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_504

module FA__2_507 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_507

module FA__2_510 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_510

module FA__2_513 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_513

module FA__2_516 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_516

module FA__2_519 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_519

module FA__2_522 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_522

module FA__2_525 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_525

module FA__2_528 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_528

module FA__2_531 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_531

module HA__2_534 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_534

module FA__2_537 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_537

module FA__2_540 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_540

module FA__2_543 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_543

module FA__2_546 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_546

module FA__2_549 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_549

module FA__2_552 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_552

module FA__2_555 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_555

module FA__2_558 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_558

module HA__2_561 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_561

module FA__2_564 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_564

module HA__2_567 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_567

module FA__2_570 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_570

module FA__2_573 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_573

module FA__2_576 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_576

module HA__2_579 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_579

module HA__2_582 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_582

module HA__2_585 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_585

module HA__2_588 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_588

module HA__2_591 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_591

module HA__2_594 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_594

module HA__2_597 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_597

module FA__2_600 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_600

module FA__2_603 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_603

module FA__2_606 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_606

module FA__2_609 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_609

module HA__2_612 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__2_612

module FA__2_615 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_615

module FA__2_618 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_618

module FA__2_621 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_621

module FA__2_624 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_624

module FA__2_627 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_627

module WTM8__2_628 (A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
wire spw_n8;
wire spw_n16;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (spw_n16));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (spw_n16));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (spw_n16));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (spw_n16));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (spw_n16));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (spw_n16));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (spw_n16));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (spw_n16));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (spw_n8));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (spw_n8));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (spw_n8));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (spw_n8));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (spw_n8));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (spw_n8));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (spw_n8));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (spw_n8));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__2_441 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__2_444 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__2_447 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__2_450 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__2_453 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__2_456 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__2_459 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__2_462 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__2_465 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__2_468 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__2_471 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__2_474 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__2_477 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__2_480 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__2_483 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__2_486 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__2_489 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__2_492 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__2_495 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__2_498 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__2_501 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__2_504 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__2_507 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__2_510 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__2_513 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__2_516 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__2_519 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__2_522 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__2_525 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__2_528 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__2_531 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__2_534 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__2_537 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__2_540 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__2_543 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__2_546 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__2_549 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__2_552 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__2_555 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__2_558 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__2_561 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__2_564 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__2_567 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__2_570 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__2_573 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__2_576 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__2_579 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__2_582 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__2_585 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__2_588 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__2_591 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__2_594 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__2_597 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__2_600 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__2_603 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__2_606 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__2_609 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__2_612 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__2_615 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__2_618 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__2_621 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__2_624 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__2_627 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));
BUF_X1 spw__L3_c7_c1 (.Z (spw_n8), .A (B[7]));
BUF_X2 spw__L3_c3_c4 (.Z (spw_n16), .A (B[5]));

endmodule //WTM8__2_628

module FA__2_1949 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1949

module FA__2_1952 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1952

module FA__2_1955 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1955

module FA__2_1958 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1958

module FA__2_1961 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1961

module FA__2_1964 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1964

module FA__2_1967 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1967

module FA__2_1970 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__2_1970

module FA__2_1973 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1973

module FA__2_1976 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1976

module FA__2_1979 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1979

module FA__2_1982 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1982

module FA__2_1985 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1985

module FA__2_1988 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1988

module FA__2_1991 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__2_1991

module FA__2_1994 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__2_1994

module adder64__2_2091 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;


FA__2_1949 genblk1_47_F (.carry (z[48]), .sum (z[47]), .b (y[47]), .cin (\carry[46] ));
FA__2_1952 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .b (y[46]), .cin (\carry[45] ));
FA__2_1955 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .b (y[45]), .cin (\carry[44] ));
FA__2_1958 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .b (y[44]), .cin (\carry[43] ));
FA__2_1961 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .b (y[43]), .cin (\carry[42] ));
FA__2_1964 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .b (y[42]), .cin (\carry[41] ));
FA__2_1967 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .b (y[41]), .cin (\carry[40] ));
FA__2_1970 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .b (y[40]), .cin (\carry[39] ));
FA__2_1973 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .a (x[39]), .b (y[39]), .cin (\carry[38] ));
FA__2_1976 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .a (x[38]), .b (y[38]), .cin (\carry[37] ));
FA__2_1979 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .a (x[37]), .b (y[37]), .cin (\carry[36] ));
FA__2_1982 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .a (x[36]), .b (y[36]), .cin (\carry[35] ));
FA__2_1985 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .a (x[35]), .b (y[35]), .cin (\carry[34] ));
FA__2_1988 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .a (x[34]), .b (y[34]), .cin (\carry[33] ));
FA__2_1991 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .a (x[33]), .b (y[33]), .cin (\carry[32] ));
FA__2_1994 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32]));

endmodule //adder64__2_2091

module FA__1_140 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_140

module HA__1_374 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_374

module FA__1_137 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_137

module FA__1_134 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_134

module HA__1_371 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_371

module FA__1_131 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_131

module FA__1_128 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_128

module HA__1_368 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_368

module FA__1_125 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_125

module FA__1_122 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_122

module FA__1_119 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_119

module HA__1_365 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_365

module FA__1_116 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_116

module HA__1_362 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_362

module FA__1_113 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_113

module FA__1_110 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_110

module FA__1_107 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_107

module FA__1_104 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_104

module FA__1_101 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_101

module FA__1_98 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_98

module FA__1_95 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_95

module FA__1_92 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_92

module FA__1_89 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_89

module FA__1_86 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_86

module FA__1_83 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_83

module FA__1_80 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_80

module FA__1_77 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_77

module FA__1_74 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_74

module FA__1_71 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_71

module FA__1_68 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_68

module FA__1_65 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_65

module HA__1_359 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_359

module FA__1_62 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_62

module FA__1_59 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_59

module FA__1_56 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_56

module FA__1_53 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_53

module FA__1_50 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_50

module FA__1_47 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_47

module FA__1_44 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_44

module FA__1_41 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_41

module HA__1_356 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_356

module FA__1_38 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_38

module HA__1_353 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_353

module FA__1_35 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_35

module FA__1_32 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_32

module FA__1_29 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_29

module HA__1_350 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_350

module HA__1_347 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_347

module HA__1_344 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_344

module HA__1_341 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_341

module HA__1_338 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_338

module HA__1_335 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_335

module HA__1_332 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_332

module FA__1_26 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_26

module FA__1_23 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_23

module FA__1_20 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_20

module FA__1_17 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_17

module HA__1_329 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_329

module FA__1_14 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_14

module FA__1_11 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_11

module FA__1_8 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_8

module FA__1_5 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_5

module FA__1_2 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2

module WTM8__0_153 (A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_140 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_374 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_137 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_134 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_371 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_131 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_128 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_368 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_125 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_122 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_119 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_365 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_116 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_362 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_113 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_110 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_107 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_104 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_101 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_98 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_95 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_92 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_89 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_86 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_83 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_80 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_77 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_74 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_71 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_68 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_65 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_359 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_62 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_59 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_56 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_53 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_50 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_47 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_44 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_41 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_356 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_38 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_353 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_35 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_32 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_29 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_350 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_347 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_344 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_341 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_338 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_335 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_332 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_26 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_23 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_20 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_17 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_329 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_14 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_11 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_8 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_5 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_2 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__0_153

module FA__0_149 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


XOR2_X1 i_0_0 (.Z (sum), .A (b), .B (cin));

endmodule //FA__0_149

module FA__1_326 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X2 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_326

module FA__1_323 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X2 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_323

module FA__1_320 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_320

module FA__1_317 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_317

module FA__1_314 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_314

module FA__1_311 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_311

module FA__1_308 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_308

module FA__1_305 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_305

module FA__1_302 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X2 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_302

module FA__1_299 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_299

module FA__1_296 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X4 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_296

module FA__1_293 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X2 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_293

module FA__1_290 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_290

module FA__1_287 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_287

module FA__1_284 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_284

module FA__1_281 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_281

module FA__1_278 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_278

module FA__1_275 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X4 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_275

module FA__1_272 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X4 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_272

module FA__1_269 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_269

module FA__1_266 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_266

module FA__1_263 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_263

module FA__1_260 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_260

module FA__1_257 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_257

module FA__1_254 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_254

module FA__1_251 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_251

module FA__1_248 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_248

module FA__1_245 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_245

module FA__1_242 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X4 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_242

module FA__1_239 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_239

module FA__1_236 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_236

module FA__1_233 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_233

module FA__1_230 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_230

module FA__1_227 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_227

module FA__1_224 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_224

module FA__1_221 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_221

module FA__1_218 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_218

module FA__1_215 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_215

module FA__1_212 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_212

module FA__1_209 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_209

module FA__1_206 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_206

module FA__1_203 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_203

module FA__1_200 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_200

module FA__1_197 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_197

module FA__1_194 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_194

module FA__1_191 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_191

module FA__1_188 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_188

module adder64__0_154 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[62] ;
wire \carry[61] ;
wire \carry[60] ;
wire \carry[59] ;
wire \carry[58] ;
wire \carry[57] ;
wire \carry[56] ;
wire \carry[55] ;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;
wire \carry[23] ;
wire \carry[22] ;
wire \carry[21] ;
wire \carry[20] ;
wire \carry[19] ;
wire \carry[18] ;
wire \carry[17] ;
wire \carry[16] ;


FA__0_149 genblk1_63_F (.sum (z[63]), .b (y[63]), .cin (\carry[62] ));
FA__1_326 genblk1_62_F (.carry (\carry[62] ), .sum (z[62]), .b (y[62]), .cin (\carry[61] ));
FA__1_323 genblk1_61_F (.carry (\carry[61] ), .sum (z[61]), .b (y[61]), .cin (\carry[60] ));
FA__1_320 genblk1_60_F (.carry (\carry[60] ), .sum (z[60]), .b (y[60]), .cin (\carry[59] ));
FA__1_317 genblk1_59_F (.carry (\carry[59] ), .sum (z[59]), .b (y[59]), .cin (\carry[58] ));
FA__1_314 genblk1_58_F (.carry (\carry[58] ), .sum (z[58]), .b (y[58]), .cin (\carry[57] ));
FA__1_311 genblk1_57_F (.carry (\carry[57] ), .sum (z[57]), .b (y[57]), .cin (\carry[56] ));
FA__1_308 genblk1_56_F (.carry (\carry[56] ), .sum (z[56]), .b (y[56]), .cin (\carry[55] ));
FA__1_305 genblk1_55_F (.carry (\carry[55] ), .sum (z[55]), .b (y[55]), .cin (\carry[54] ));
FA__1_302 genblk1_54_F (.carry (\carry[54] ), .sum (z[54]), .b (y[54]), .cin (\carry[53] ));
FA__1_299 genblk1_53_F (.carry (\carry[53] ), .sum (z[53]), .b (y[53]), .cin (\carry[52] ));
FA__1_296 genblk1_52_F (.carry (\carry[52] ), .sum (z[52]), .b (y[52]), .cin (\carry[51] ));
FA__1_293 genblk1_51_F (.carry (\carry[51] ), .sum (z[51]), .b (y[51]), .cin (\carry[50] ));
FA__1_290 genblk1_50_F (.carry (\carry[50] ), .sum (z[50]), .a (x[50]), .b (y[50]), .cin (\carry[49] ));
FA__1_287 genblk1_49_F (.carry (\carry[49] ), .sum (z[49]), .a (x[49]), .b (y[49])
    , .cin (\carry[48] ));
FA__1_284 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .a (x[48]), .b (y[48]), .cin (\carry[47] ));
FA__1_281 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .a (x[47]), .b (y[47])
    , .cin (\carry[46] ));
FA__1_278 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .a (x[46]), .b (y[46]), .cin (\carry[45] ));
FA__1_275 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .a (x[45]), .b (y[45]), .cin (\carry[44] ));
FA__1_272 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .a (x[44]), .b (y[44]), .cin (\carry[43] ));
FA__1_269 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .a (x[43]), .b (y[43]), .cin (\carry[42] ));
FA__1_266 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .a (x[42]), .b (y[42])
    , .cin (\carry[41] ));
FA__1_263 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .a (x[41]), .b (y[41])
    , .cin (\carry[40] ));
FA__1_260 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .a (x[40]), .b (y[40])
    , .cin (\carry[39] ));
FA__1_257 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .a (x[39]), .b (y[39])
    , .cin (\carry[38] ));
FA__1_254 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .a (x[38]), .b (y[38])
    , .cin (\carry[37] ));
FA__1_251 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .a (x[37]), .b (y[37])
    , .cin (\carry[36] ));
FA__1_248 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .a (x[36]), .b (y[36])
    , .cin (\carry[35] ));
FA__1_245 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .a (x[35]), .b (y[35])
    , .cin (\carry[34] ));
FA__1_242 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .a (x[34]), .b (y[34]), .cin (\carry[33] ));
FA__1_239 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .a (x[33]), .b (y[33])
    , .cin (\carry[32] ));
FA__1_236 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32])
    , .cin (\carry[31] ));
FA__1_233 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .a (x[31]), .b (y[31])
    , .cin (\carry[30] ));
FA__1_230 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .a (x[30]), .b (y[30])
    , .cin (\carry[29] ));
FA__1_227 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .a (x[29]), .b (y[29]), .cin (\carry[28] ));
FA__1_224 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .a (x[28]), .b (y[28])
    , .cin (\carry[27] ));
FA__1_221 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .a (x[27]), .b (y[27]), .cin (\carry[26] ));
FA__1_218 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .a (x[26]), .b (y[26])
    , .cin (\carry[25] ));
FA__1_215 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .a (x[25]), .b (y[25])
    , .cin (\carry[24] ));
FA__1_212 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24])
    , .cin (\carry[23] ));
FA__1_209 genblk1_23_F (.carry (\carry[23] ), .sum (z[23]), .a (x[23]), .b (y[23])
    , .cin (\carry[22] ));
FA__1_206 genblk1_22_F (.carry (\carry[22] ), .sum (z[22]), .a (x[22]), .b (y[22])
    , .cin (\carry[21] ));
FA__1_203 genblk1_21_F (.carry (\carry[21] ), .sum (z[21]), .a (x[21]), .b (y[21])
    , .cin (\carry[20] ));
FA__1_200 genblk1_20_F (.carry (\carry[20] ), .sum (z[20]), .a (x[20]), .b (y[20])
    , .cin (\carry[19] ));
FA__1_197 genblk1_19_F (.carry (\carry[19] ), .sum (z[19]), .a (x[19]), .b (y[19])
    , .cin (\carry[18] ));
FA__1_194 genblk1_18_F (.carry (\carry[18] ), .sum (z[18]), .a (x[18]), .b (y[18])
    , .cin (\carry[17] ));
FA__1_191 genblk1_17_F (.carry (\carry[17] ), .sum (z[17]), .a (x[17]), .b (y[17])
    , .cin (\carry[16] ));
FA__1_188 genblk1_16_F (.carry (\carry[16] ), .sum (z[16]), .a (x[16]), .b (y[16]));

endmodule //adder64__0_154

module datapath (p_0, out);

output [63:0] p_0;
input [63:0] out;
wire n_61;
wire n_0;
wire n_60;
wire n_59;
wire n_58;
wire n_1;
wire n_57;
wire n_56;
wire n_2;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_3;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_4;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_5;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;


INV_X1 i_135 (.ZN (n_72), .A (out[60]));
INV_X1 i_134 (.ZN (n_71), .A (out[55]));
INV_X1 i_133 (.ZN (n_70), .A (out[51]));
INV_X1 i_132 (.ZN (n_69), .A (out[42]));
INV_X1 i_131 (.ZN (n_68), .A (out[40]));
INV_X1 i_130 (.ZN (n_67), .A (out[36]));
INV_X1 i_129 (.ZN (n_66), .A (out[31]));
INV_X1 i_128 (.ZN (n_65), .A (out[26]));
INV_X1 i_127 (.ZN (n_64), .A (out[21]));
INV_X1 i_126 (.ZN (n_63), .A (out[13]));
INV_X1 i_125 (.ZN (n_62), .A (out[11]));
OR3_X1 i_124 (.ZN (n_61), .A1 (out[2]), .A2 (out[1]), .A3 (out[0]));
OR2_X1 i_123 (.ZN (n_60), .A1 (n_61), .A2 (out[3]));
OR2_X1 i_122 (.ZN (n_59), .A1 (n_60), .A2 (out[4]));
OR3_X1 i_121 (.ZN (n_58), .A1 (n_59), .A2 (out[5]), .A3 (out[6]));
OR2_X1 i_120 (.ZN (n_57), .A1 (n_58), .A2 (out[7]));
OR3_X1 i_119 (.ZN (n_56), .A1 (n_57), .A2 (out[8]), .A3 (out[9]));
NOR2_X1 i_118 (.ZN (n_55), .A1 (n_56), .A2 (out[10]));
NAND2_X1 i_117 (.ZN (n_54), .A1 (n_55), .A2 (n_62));
NOR2_X1 i_116 (.ZN (n_53), .A1 (n_54), .A2 (out[12]));
NAND2_X1 i_115 (.ZN (n_52), .A1 (n_53), .A2 (n_63));
OR3_X1 i_114 (.ZN (n_51), .A1 (n_52), .A2 (out[14]), .A3 (out[15]));
OR2_X1 i_113 (.ZN (n_50), .A1 (n_51), .A2 (out[16]));
OR2_X1 i_112 (.ZN (n_49), .A1 (n_50), .A2 (out[17]));
NOR2_X1 i_111 (.ZN (n_48), .A1 (n_49), .A2 (out[18]));
NOR3_X1 i_110 (.ZN (n_47), .A1 (n_49), .A2 (out[18]), .A3 (out[19]));
NOR4_X1 i_109 (.ZN (n_46), .A1 (n_49), .A2 (out[18]), .A3 (out[19]), .A4 (out[20]));
NAND2_X1 i_108 (.ZN (n_45), .A1 (n_46), .A2 (n_64));
OR2_X1 i_107 (.ZN (n_44), .A1 (n_45), .A2 (out[22]));
NOR2_X1 i_106 (.ZN (n_43), .A1 (n_44), .A2 (out[23]));
NOR3_X1 i_105 (.ZN (n_42), .A1 (n_44), .A2 (out[23]), .A3 (out[24]));
NOR4_X1 i_104 (.ZN (n_41), .A1 (n_44), .A2 (out[23]), .A3 (out[24]), .A4 (out[25]));
NAND2_X1 i_103 (.ZN (n_40), .A1 (n_41), .A2 (n_65));
OR2_X1 i_102 (.ZN (n_39), .A1 (n_40), .A2 (out[27]));
NOR2_X1 i_101 (.ZN (n_38), .A1 (n_39), .A2 (out[28]));
NOR3_X1 i_100 (.ZN (n_37), .A1 (n_39), .A2 (out[28]), .A3 (out[29]));
NOR4_X1 i_99 (.ZN (n_36), .A1 (n_39), .A2 (out[28]), .A3 (out[29]), .A4 (out[30]));
NAND2_X1 i_98 (.ZN (n_35), .A1 (n_36), .A2 (n_66));
OR2_X1 i_97 (.ZN (n_34), .A1 (n_35), .A2 (out[32]));
NOR2_X1 i_96 (.ZN (n_33), .A1 (n_34), .A2 (out[33]));
NOR3_X1 i_95 (.ZN (n_32), .A1 (n_34), .A2 (out[33]), .A3 (out[34]));
NOR4_X1 i_94 (.ZN (n_31), .A1 (n_34), .A2 (out[33]), .A3 (out[34]), .A4 (out[35]));
NAND2_X1 i_93 (.ZN (n_30), .A1 (n_31), .A2 (n_67));
OR2_X1 i_92 (.ZN (n_29), .A1 (n_30), .A2 (out[37]));
NOR2_X1 i_91 (.ZN (n_28), .A1 (n_29), .A2 (out[38]));
NOR3_X1 i_90 (.ZN (n_27), .A1 (n_29), .A2 (out[38]), .A3 (out[39]));
NAND2_X1 i_89 (.ZN (n_26), .A1 (n_27), .A2 (n_68));
NOR2_X1 i_88 (.ZN (n_25), .A1 (n_26), .A2 (out[41]));
NAND2_X1 i_87 (.ZN (n_24), .A1 (n_25), .A2 (n_69));
OR3_X1 i_86 (.ZN (n_23), .A1 (n_24), .A2 (out[43]), .A3 (out[44]));
OR2_X1 i_85 (.ZN (n_22), .A1 (n_23), .A2 (out[45]));
OR2_X1 i_84 (.ZN (n_21), .A1 (n_22), .A2 (out[46]));
OR2_X1 i_83 (.ZN (n_20), .A1 (n_21), .A2 (out[47]));
NOR2_X1 i_82 (.ZN (n_19), .A1 (n_20), .A2 (out[48]));
NOR3_X1 i_81 (.ZN (n_18), .A1 (n_20), .A2 (out[48]), .A3 (out[49]));
NOR4_X4 i_80 (.ZN (n_17), .A1 (n_20), .A2 (out[48]), .A3 (out[49]), .A4 (out[50]));
NAND2_X4 i_79 (.ZN (n_16), .A1 (n_17), .A2 (n_70));
NOR2_X1 i_78 (.ZN (n_15), .A1 (n_16), .A2 (out[52]));
NOR3_X1 i_77 (.ZN (n_14), .A1 (n_16), .A2 (out[52]), .A3 (out[53]));
NOR4_X4 i_76 (.ZN (n_13), .A1 (n_16), .A2 (out[52]), .A3 (out[53]), .A4 (out[54]));
NAND2_X2 i_75 (.ZN (n_12), .A1 (n_13), .A2 (n_71));
OR3_X4 i_74 (.ZN (n_11), .A1 (n_12), .A2 (out[56]), .A3 (out[57]));
NOR2_X1 i_73 (.ZN (n_10), .A1 (n_11), .A2 (out[58]));
NOR3_X4 i_72 (.ZN (n_9), .A1 (n_11), .A2 (out[58]), .A3 (out[59]));
NAND2_X4 i_71 (.ZN (n_8), .A1 (n_9), .A2 (n_72));
NOR2_X1 i_70 (.ZN (n_7), .A1 (n_8), .A2 (out[61]));
NOR3_X4 i_69 (.ZN (n_6), .A1 (n_8), .A2 (out[61]), .A3 (out[62]));
XNOR2_X1 i_68 (.ZN (p_0[63]), .A (out[63]), .B (n_6));
XNOR2_X1 i_67 (.ZN (p_0[62]), .A (out[62]), .B (n_7));
XOR2_X1 i_66 (.Z (p_0[61]), .A (out[61]), .B (n_8));
XNOR2_X1 i_65 (.ZN (p_0[60]), .A (out[60]), .B (n_9));
XNOR2_X1 i_64 (.ZN (p_0[59]), .A (out[59]), .B (n_10));
XOR2_X1 i_63 (.Z (p_0[58]), .A (out[58]), .B (n_11));
OAI21_X1 i_62 (.ZN (n_5), .A (out[57]), .B1 (n_12), .B2 (out[56]));
AND2_X2 i_61 (.ZN (p_0[57]), .A1 (n_11), .A2 (n_5));
XOR2_X1 i_60 (.Z (p_0[56]), .A (out[56]), .B (n_12));
XNOR2_X1 i_59 (.ZN (p_0[55]), .A (out[55]), .B (n_13));
XNOR2_X1 i_58 (.ZN (p_0[54]), .A (out[54]), .B (n_14));
XNOR2_X1 i_57 (.ZN (p_0[53]), .A (out[53]), .B (n_15));
XOR2_X1 i_56 (.Z (p_0[52]), .A (out[52]), .B (n_16));
XNOR2_X1 i_55 (.ZN (p_0[51]), .A (out[51]), .B (n_17));
XNOR2_X1 i_54 (.ZN (p_0[50]), .A (out[50]), .B (n_18));
XNOR2_X1 i_53 (.ZN (p_0[49]), .A (out[49]), .B (n_19));
XOR2_X1 i_52 (.Z (p_0[48]), .A (out[48]), .B (n_20));
XOR2_X1 i_51 (.Z (p_0[47]), .A (out[47]), .B (n_21));
XOR2_X1 i_50 (.Z (p_0[46]), .A (out[46]), .B (n_22));
XOR2_X1 i_49 (.Z (p_0[45]), .A (out[45]), .B (n_23));
OAI21_X1 i_48 (.ZN (n_4), .A (out[44]), .B1 (n_24), .B2 (out[43]));
AND2_X1 i_47 (.ZN (p_0[44]), .A1 (n_23), .A2 (n_4));
XOR2_X1 i_46 (.Z (p_0[43]), .A (out[43]), .B (n_24));
XNOR2_X1 i_45 (.ZN (p_0[42]), .A (out[42]), .B (n_25));
XOR2_X1 i_44 (.Z (p_0[41]), .A (out[41]), .B (n_26));
XNOR2_X1 i_43 (.ZN (p_0[40]), .A (out[40]), .B (n_27));
XNOR2_X1 i_42 (.ZN (p_0[39]), .A (out[39]), .B (n_28));
XOR2_X1 i_41 (.Z (p_0[38]), .A (out[38]), .B (n_29));
XOR2_X1 i_40 (.Z (p_0[37]), .A (out[37]), .B (n_30));
XNOR2_X1 i_39 (.ZN (p_0[36]), .A (out[36]), .B (n_31));
XNOR2_X1 i_38 (.ZN (p_0[35]), .A (out[35]), .B (n_32));
XNOR2_X1 i_37 (.ZN (p_0[34]), .A (out[34]), .B (n_33));
XOR2_X1 i_36 (.Z (p_0[33]), .A (out[33]), .B (n_34));
XOR2_X1 i_35 (.Z (p_0[32]), .A (out[32]), .B (n_35));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (out[31]), .B (n_36));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (out[30]), .B (n_37));
XNOR2_X1 i_32 (.ZN (p_0[29]), .A (out[29]), .B (n_38));
XOR2_X1 i_31 (.Z (p_0[28]), .A (out[28]), .B (n_39));
XOR2_X1 i_30 (.Z (p_0[27]), .A (out[27]), .B (n_40));
XNOR2_X1 i_29 (.ZN (p_0[26]), .A (out[26]), .B (n_41));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (out[25]), .B (n_42));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (out[24]), .B (n_43));
XOR2_X1 i_26 (.Z (p_0[23]), .A (out[23]), .B (n_44));
XOR2_X1 i_25 (.Z (p_0[22]), .A (out[22]), .B (n_45));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (out[21]), .B (n_46));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (out[20]), .B (n_47));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (out[19]), .B (n_48));
XOR2_X1 i_21 (.Z (p_0[18]), .A (out[18]), .B (n_49));
XOR2_X1 i_20 (.Z (p_0[17]), .A (out[17]), .B (n_50));
XOR2_X1 i_19 (.Z (p_0[16]), .A (out[16]), .B (n_51));
OAI21_X1 i_18 (.ZN (n_3), .A (out[15]), .B1 (n_52), .B2 (out[14]));
AND2_X1 i_17 (.ZN (p_0[15]), .A1 (n_51), .A2 (n_3));
XOR2_X1 i_16 (.Z (p_0[14]), .A (out[14]), .B (n_52));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (out[13]), .B (n_53));
XOR2_X1 i_14 (.Z (p_0[12]), .A (out[12]), .B (n_54));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (out[11]), .B (n_55));
XOR2_X1 i_12 (.Z (p_0[10]), .A (out[10]), .B (n_56));
OAI21_X1 i_11 (.ZN (n_2), .A (out[9]), .B1 (n_57), .B2 (out[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_56), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (out[8]), .B (n_57));
XOR2_X1 i_8 (.Z (p_0[7]), .A (out[7]), .B (n_58));
OAI21_X1 i_7 (.ZN (n_1), .A (out[6]), .B1 (n_59), .B2 (out[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_58), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (out[5]), .B (n_59));
XOR2_X1 i_4 (.Z (p_0[4]), .A (out[4]), .B (n_60));
XOR2_X1 i_3 (.Z (p_0[3]), .A (out[3]), .B (n_61));
OAI21_X1 i_2 (.ZN (n_0), .A (out[2]), .B1 (out[1]), .B2 (out[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_61), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (out[1]), .B (out[0]));

endmodule //datapath

module FA__1_2219 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_2219

module HA__1_2222 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2222

module FA__1_2225 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2225

module FA__1_2228 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2228

module HA__1_2231 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2231

module FA__1_2234 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2234

module FA__1_2237 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2237

module HA__1_2240 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2240

module FA__1_2243 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2243

module FA__1_2246 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2246

module FA__1_2249 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2249

module HA__1_2252 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2252

module FA__1_2255 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2255

module HA__1_2258 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2258

module FA__1_2261 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2261

module FA__1_2264 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2264

module FA__1_2267 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2267

module FA__1_2270 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2270

module FA__1_2273 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2273

module FA__1_2276 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2276

module FA__1_2279 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2279

module FA__1_2282 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2282

module FA__1_2285 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2285

module FA__1_2288 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2288

module FA__1_2291 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2291

module FA__1_2294 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2294

module FA__1_2297 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2297

module FA__1_2300 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2300

module FA__1_2303 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2303

module FA__1_2306 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2306

module FA__1_2309 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2309

module HA__1_2312 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2312

module FA__1_2315 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2315

module FA__1_2318 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2318

module FA__1_2321 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2321

module FA__1_2324 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2324

module FA__1_2327 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2327

module FA__1_2330 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2330

module FA__1_2333 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2333

module FA__1_2336 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2336

module HA__1_2339 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2339

module FA__1_2342 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2342

module HA__1_2345 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2345

module FA__1_2348 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2348

module FA__1_2351 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2351

module FA__1_2354 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2354

module HA__1_2357 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2357

module HA__1_2360 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2360

module HA__1_2363 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2363

module HA__1_2366 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2366

module HA__1_2369 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2369

module HA__1_2372 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2372

module HA__1_2375 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2375

module FA__1_2378 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2378

module FA__1_2381 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2381

module FA__1_2384 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2384

module FA__1_2387 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2387

module HA__1_2390 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2390

module FA__1_2393 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2393

module FA__1_2396 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2396

module FA__1_2399 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2399

module FA__1_2402 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2402

module FA__1_2405 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2405

module WTM8__1_2406 (A_5_PP_0, A_5_PP_1, A_3_PP_0, A_4_PP_0, A_4_PP_1, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_5_PP_0;
input A_5_PP_1;
input A_3_PP_0;
input A_4_PP_0;
input A_4_PP_1;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A_4_PP_1), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A_3_PP_0), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A_5_PP_1), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A_3_PP_0), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A_5_PP_1), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A_4_PP_0), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A_5_PP_0), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A_4_PP_0), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A_3_PP_0), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A_5_PP_0), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A_4_PP_0), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A_3_PP_0), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A_5_PP_0), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A_3_PP_0), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A_5_PP_0), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A_3_PP_0), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_2219 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_2222 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_2225 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_2228 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_2231 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_2234 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_2237 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_2240 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_2243 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_2246 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_2249 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_2252 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_2255 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_2258 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_2261 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_2264 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_2267 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_2270 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_2273 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_2276 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_2279 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_2282 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_2285 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_2288 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_2291 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_2294 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_2297 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_2300 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_2303 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_2306 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_2309 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_2312 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_2315 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_2318 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_2321 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_2324 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_2327 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_2330 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_2333 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_2336 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_2339 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_2342 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_2345 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_2348 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_2351 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_2354 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_2357 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_2360 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_2363 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_2366 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_2369 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_2372 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_2375 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_2378 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_2381 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_2384 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_2387 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_2390 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_2393 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_2396 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_2399 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_2402 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_2405 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__1_2406

module datapath__0_79 (p_0, A);

output [31:0] p_0;
input [31:0] A;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (A[25]));
INV_X1 i_63 (.ZN (n_32), .A (A[21]));
INV_X1 i_62 (.ZN (n_31), .A (A[14]));
INV_X1 i_61 (.ZN (n_30), .A (A[11]));
OR3_X4 i_60 (.ZN (n_29), .A1 (A[2]), .A2 (A[1]), .A3 (A[0]));
OR2_X4 i_59 (.ZN (n_28), .A1 (n_29), .A2 (A[3]));
OR2_X4 i_58 (.ZN (n_27), .A1 (n_28), .A2 (A[4]));
OR3_X4 i_57 (.ZN (n_26), .A1 (n_27), .A2 (A[5]), .A3 (A[6]));
OR2_X2 i_56 (.ZN (n_25), .A1 (n_26), .A2 (A[7]));
OR3_X4 i_55 (.ZN (n_24), .A1 (n_25), .A2 (A[8]), .A3 (A[9]));
NOR2_X4 i_54 (.ZN (n_23), .A1 (n_24), .A2 (A[10]));
NAND2_X2 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (A[12]));
NOR3_X4 i_51 (.ZN (n_20), .A1 (n_22), .A2 (A[12]), .A3 (A[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (A[15]), .A3 (A[16]));
OR2_X4 i_48 (.ZN (n_17), .A1 (n_18), .A2 (A[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (A[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (A[18]), .A3 (A[19]));
NOR4_X4 i_45 (.ZN (n_14), .A1 (n_17), .A2 (A[18]), .A3 (A[19]), .A4 (A[20]));
NAND2_X2 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (A[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (A[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (A[23]), .A3 (A[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (A[26]), .A3 (A[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (A[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (A[28]), .A3 (A[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (A[28]), .A3 (A[29]), .A4 (A[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (A[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (A[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (A[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (A[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (A[27]), .B1 (n_9), .B2 (A[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (A[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (A[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (A[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (A[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (A[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (A[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (A[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (A[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (A[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (A[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (A[16]), .B1 (n_19), .B2 (A[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (A[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (A[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (A[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (A[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (A[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (A[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (A[9]), .B1 (n_25), .B2 (A[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (A[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (A[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (A[6]), .B1 (n_27), .B2 (A[5]));
AND2_X2 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (A[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (A[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (A[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (A[2]), .B1 (A[1]), .B2 (A[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (A[1]), .B (A[0]));

endmodule //datapath__0_79

module datapath__0_81 (p_0, B);

output [31:0] p_0;
input [31:0] B;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (B[25]));
INV_X1 i_63 (.ZN (n_32), .A (B[21]));
INV_X1 i_62 (.ZN (n_31), .A (B[14]));
INV_X1 i_61 (.ZN (n_30), .A (B[11]));
OR3_X4 i_60 (.ZN (n_29), .A1 (B[2]), .A2 (B[1]), .A3 (B[0]));
OR2_X4 i_59 (.ZN (n_28), .A1 (n_29), .A2 (B[3]));
OR2_X2 i_58 (.ZN (n_27), .A1 (n_28), .A2 (B[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (B[5]), .A3 (B[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (B[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (B[8]), .A3 (B[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (B[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (B[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (B[12]), .A3 (B[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (B[15]), .A3 (B[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (B[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (B[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (B[18]), .A3 (B[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (B[18]), .A3 (B[19]), .A4 (B[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (B[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (B[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (B[23]), .A3 (B[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (B[26]), .A3 (B[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (B[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (B[28]), .A3 (B[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (B[28]), .A3 (B[29]), .A4 (B[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (B[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (B[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (B[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (B[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (B[27]), .B1 (n_9), .B2 (B[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (B[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (B[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (B[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (B[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (B[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (B[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (B[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (B[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (B[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (B[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (B[16]), .B1 (n_19), .B2 (B[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (B[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (B[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (B[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (B[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (B[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (B[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (B[9]), .B1 (n_25), .B2 (B[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (B[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (B[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (B[6]), .B1 (n_27), .B2 (B[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (B[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (B[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (B[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (B[2]), .B1 (B[1]), .B2 (B[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (B[1]), .B (B[0]));

endmodule //datapath__0_81

module FA__1_3609 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3609

module FA__1_3612 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3612

module FA__1_3615 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3615

module FA__1_3618 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3618

module FA__1_3621 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3621

module FA__1_3624 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3624

module FA__1_3627 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3627

module FA__1_3630 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3630

module FA__1_3633 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3633

module FA__1_3636 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3636

module FA__1_3639 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3639

module FA__1_3642 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3642

module FA__1_3645 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3645

module FA__1_3648 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3648

module FA__1_3651 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3651

module FA__1_3654 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3654

module FA__1_3657 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3657

module FA__1_3660 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3660

module FA__1_3663 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3663

module FA__1_3666 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3666

module FA__1_3669 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3669

module FA__1_3672 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3672

module FA__1_3675 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3675

module FA__1_3678 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3678

module FA__1_3681 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3681

module FA__1_3684 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3684

module FA__1_3687 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3687

module FA__1_3690 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3690

module FA__1_3693 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3693

module FA__1_3696 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3696

module FA__1_3699 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3699

module FA__1_3702 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3702

module FA__1_3705 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3705

module FA__1_3708 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3708

module FA__1_3711 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3711

module FA__1_3714 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3714

module FA__1_3717 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3717

module FA__1_3720 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3720

module FA__1_3723 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3723

module FA__1_3726 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3726

module FA__1_3729 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3729

module FA__1_3732 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_3732

module adder64__1_3757 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;
wire \carry[23] ;
wire \carry[22] ;
wire \carry[21] ;
wire \carry[20] ;
wire \carry[19] ;
wire \carry[18] ;
wire \carry[17] ;
wire \carry[16] ;
wire \carry[15] ;
wire \carry[14] ;
wire \carry[13] ;
wire \carry[12] ;
wire \carry[11] ;
wire \carry[10] ;
wire \carry[9] ;
wire \carry[8] ;


FA__1_3609 genblk1_49_F (.carry (z[50]), .sum (z[49]), .b (y[49]), .cin (\carry[48] ));
FA__1_3612 genblk1_48_F (.carry (\carry[48] ), .sum (z[48]), .b (y[48]), .cin (\carry[47] ));
FA__1_3615 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .b (y[47]), .cin (\carry[46] ));
FA__1_3618 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .b (y[46]), .cin (\carry[45] ));
FA__1_3621 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .b (y[45]), .cin (\carry[44] ));
FA__1_3624 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .b (y[44]), .cin (\carry[43] ));
FA__1_3627 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .b (y[43]), .cin (\carry[42] ));
FA__1_3630 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .b (y[42]), .cin (\carry[41] ));
FA__1_3633 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .a (x[41]), .b (y[41]), .cin (\carry[40] ));
FA__1_3636 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .a (x[40]), .b (y[40]), .cin (\carry[39] ));
FA__1_3639 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .a (x[39]), .b (y[39]), .cin (\carry[38] ));
FA__1_3642 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .a (x[38]), .b (y[38]), .cin (\carry[37] ));
FA__1_3645 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .a (x[37]), .b (y[37])
    , .cin (\carry[36] ));
FA__1_3648 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .a (x[36]), .b (y[36])
    , .cin (\carry[35] ));
FA__1_3651 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .a (x[35]), .b (y[35]), .cin (\carry[34] ));
FA__1_3654 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .a (x[34]), .b (y[34])
    , .cin (\carry[33] ));
FA__1_3657 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .a (x[33]), .b (y[33])
    , .cin (\carry[32] ));
FA__1_3660 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32])
    , .cin (\carry[31] ));
FA__1_3663 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .a (x[31]), .b (y[31])
    , .cin (\carry[30] ));
FA__1_3666 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .a (x[30]), .b (y[30])
    , .cin (\carry[29] ));
FA__1_3669 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .a (x[29]), .b (y[29]), .cin (\carry[28] ));
FA__1_3672 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .a (x[28]), .b (y[28])
    , .cin (\carry[27] ));
FA__1_3675 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .a (x[27]), .b (y[27])
    , .cin (\carry[26] ));
FA__1_3678 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .a (x[26]), .b (y[26])
    , .cin (\carry[25] ));
FA__1_3681 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .a (x[25]), .b (y[25])
    , .cin (\carry[24] ));
FA__1_3684 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24])
    , .cin (\carry[23] ));
FA__1_3687 genblk1_23_F (.carry (\carry[23] ), .sum (z[23]), .a (x[23]), .b (y[23])
    , .cin (\carry[22] ));
FA__1_3690 genblk1_22_F (.carry (\carry[22] ), .sum (z[22]), .a (x[22]), .b (y[22]), .cin (\carry[21] ));
FA__1_3693 genblk1_21_F (.carry (\carry[21] ), .sum (z[21]), .a (x[21]), .b (y[21])
    , .cin (\carry[20] ));
FA__1_3696 genblk1_20_F (.carry (\carry[20] ), .sum (z[20]), .a (x[20]), .b (y[20])
    , .cin (\carry[19] ));
FA__1_3699 genblk1_19_F (.carry (\carry[19] ), .sum (z[19]), .a (x[19]), .b (y[19]), .cin (\carry[18] ));
FA__1_3702 genblk1_18_F (.carry (\carry[18] ), .sum (z[18]), .a (x[18]), .b (y[18])
    , .cin (\carry[17] ));
FA__1_3705 genblk1_17_F (.carry (\carry[17] ), .sum (z[17]), .a (x[17]), .b (y[17]), .cin (\carry[16] ));
FA__1_3708 genblk1_16_F (.carry (\carry[16] ), .sum (z[16]), .a (x[16]), .b (y[16])
    , .cin (\carry[15] ));
FA__1_3711 genblk1_15_F (.carry (\carry[15] ), .sum (z[15]), .a (x[15]), .b (y[15])
    , .cin (\carry[14] ));
FA__1_3714 genblk1_14_F (.carry (\carry[14] ), .sum (z[14]), .a (x[14]), .b (y[14])
    , .cin (\carry[13] ));
FA__1_3717 genblk1_13_F (.carry (\carry[13] ), .sum (z[13]), .a (x[13]), .b (y[13])
    , .cin (\carry[12] ));
FA__1_3720 genblk1_12_F (.carry (\carry[12] ), .sum (z[12]), .a (x[12]), .b (y[12])
    , .cin (\carry[11] ));
FA__1_3723 genblk1_11_F (.carry (\carry[11] ), .sum (z[11]), .a (x[11]), .b (y[11])
    , .cin (\carry[10] ));
FA__1_3726 genblk1_10_F (.carry (\carry[10] ), .sum (z[10]), .a (x[10]), .b (y[10])
    , .cin (\carry[9] ));
FA__1_3729 genblk1_9_F (.carry (\carry[9] ), .sum (z[9]), .a (x[9]), .b (y[9]), .cin (\carry[8] ));
FA__1_3732 genblk1_8_F (.carry (\carry[8] ), .sum (z[8]), .a (x[8]), .b (y[8]));

endmodule //adder64__1_3757

module FA__1_3419 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3419

module FA__1_3422 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3422

module FA__1_3425 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3425

module FA__1_3428 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3428

module FA__1_3431 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3431

module FA__1_3434 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3434

module FA__1_3437 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3437

module FA__1_3440 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3440

module FA__1_3443 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3443

module FA__1_3446 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3446

module FA__1_3449 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3449

module FA__1_3452 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3452

module FA__1_3455 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3455

module FA__1_3458 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3458

module FA__1_3461 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3461

module FA__1_3464 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3464

module FA__1_3467 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3467

module FA__1_3470 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3470

module FA__1_3473 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3473

module FA__1_3476 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3476

module FA__1_3479 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3479

module FA__1_3482 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3482

module FA__1_3485 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3485

module FA__1_3488 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3488

module FA__1_3491 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_3491

module adder64__1_3564 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;


FA__1_3419 genblk1_48_F (.carry (z[49]), .sum (z[48]), .b (y[48]), .cin (\carry[47] ));
FA__1_3422 genblk1_47_F (.carry (\carry[47] ), .sum (z[47]), .b (y[47]), .cin (\carry[46] ));
FA__1_3425 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .b (y[46]), .cin (\carry[45] ));
FA__1_3428 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .b (y[45]), .cin (\carry[44] ));
FA__1_3431 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .b (y[44]), .cin (\carry[43] ));
FA__1_3434 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .b (y[43]), .cin (\carry[42] ));
FA__1_3437 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .b (y[42]), .cin (\carry[41] ));
FA__1_3440 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .b (y[41]), .cin (\carry[40] ));
FA__1_3443 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .b (y[40]), .cin (\carry[39] ));
FA__1_3446 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .b (y[39]), .cin (\carry[38] ));
FA__1_3449 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .b (y[38]), .cin (\carry[37] ));
FA__1_3452 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .b (y[37]), .cin (\carry[36] ));
FA__1_3455 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .b (y[36]), .cin (\carry[35] ));
FA__1_3458 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .b (y[35]), .cin (\carry[34] ));
FA__1_3461 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .b (y[34]), .cin (\carry[33] ));
FA__1_3464 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .b (y[33]), .cin (\carry[32] ));
FA__1_3467 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32]), .cin (\carry[31] ));
FA__1_3470 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .a (x[31]), .b (y[31]), .cin (\carry[30] ));
FA__1_3473 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .a (x[30]), .b (y[30]), .cin (\carry[29] ));
FA__1_3476 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .a (x[29]), .b (y[29]), .cin (\carry[28] ));
FA__1_3479 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .a (x[28]), .b (y[28]), .cin (\carry[27] ));
FA__1_3482 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .a (x[27]), .b (y[27]), .cin (\carry[26] ));
FA__1_3485 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .a (x[26]), .b (y[26]), .cin (\carry[25] ));
FA__1_3488 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .a (x[25]), .b (y[25]), .cin (\carry[24] ));
FA__1_3491 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24]));

endmodule //adder64__1_3564

module FA__1_3229 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3229

module FA__1_3232 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3232

module FA__1_3235 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3235

module FA__1_3238 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3238

module FA__1_3241 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3241

module FA__1_3244 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3244

module FA__1_3247 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3247

module FA__1_3250 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3250

module FA__1_3253 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3253

module FA__1_3256 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3256

module FA__1_3259 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3259

module FA__1_3262 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3262

module FA__1_3265 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3265

module FA__1_3268 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3268

module FA__1_3271 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3271

module FA__1_3274 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_3274

module adder64__1_3371 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;


FA__1_3229 genblk1_47_F (.carry (z[48]), .sum (z[47]), .b (y[47]), .cin (\carry[46] ));
FA__1_3232 genblk1_46_F (.carry (\carry[46] ), .sum (z[46]), .b (y[46]), .cin (\carry[45] ));
FA__1_3235 genblk1_45_F (.carry (\carry[45] ), .sum (z[45]), .b (y[45]), .cin (\carry[44] ));
FA__1_3238 genblk1_44_F (.carry (\carry[44] ), .sum (z[44]), .b (y[44]), .cin (\carry[43] ));
FA__1_3241 genblk1_43_F (.carry (\carry[43] ), .sum (z[43]), .b (y[43]), .cin (\carry[42] ));
FA__1_3244 genblk1_42_F (.carry (\carry[42] ), .sum (z[42]), .b (y[42]), .cin (\carry[41] ));
FA__1_3247 genblk1_41_F (.carry (\carry[41] ), .sum (z[41]), .b (y[41]), .cin (\carry[40] ));
FA__1_3250 genblk1_40_F (.carry (\carry[40] ), .sum (z[40]), .b (y[40]), .cin (\carry[39] ));
FA__1_3253 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .a (x[39]), .b (y[39]), .cin (\carry[38] ));
FA__1_3256 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .a (x[38]), .b (y[38]), .cin (\carry[37] ));
FA__1_3259 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .a (x[37]), .b (y[37]), .cin (\carry[36] ));
FA__1_3262 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .a (x[36]), .b (y[36]), .cin (\carry[35] ));
FA__1_3265 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .a (x[35]), .b (y[35]), .cin (\carry[34] ));
FA__1_3268 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .a (x[34]), .b (y[34]), .cin (\carry[33] ));
FA__1_3271 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .a (x[33]), .b (y[33]), .cin (\carry[32] ));
FA__1_3274 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .a (x[32]), .b (y[32]));

endmodule //adder64__1_3371

module FA__1_1965 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_1965

module HA__1_1968 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1968

module FA__1_1971 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1971

module FA__1_1974 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1974

module HA__1_1977 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1977

module FA__1_1980 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1980

module FA__1_1983 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1983

module HA__1_1986 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1986

module FA__1_1989 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1989

module FA__1_1992 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1992

module FA__1_1995 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1995

module HA__1_1998 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1998

module FA__1_2001 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2001

module HA__1_2004 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2004

module FA__1_2007 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2007

module FA__1_2010 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2010

module FA__1_2013 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2013

module FA__1_2016 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2016

module FA__1_2019 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2019

module FA__1_2022 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2022

module FA__1_2025 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2025

module FA__1_2028 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2028

module FA__1_2031 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2031

module FA__1_2034 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2034

module FA__1_2037 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2037

module FA__1_2040 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2040

module FA__1_2043 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2043

module FA__1_2046 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2046

module FA__1_2049 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2049

module FA__1_2052 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2052

module FA__1_2055 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2055

module HA__1_2058 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2058

module FA__1_2061 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2061

module FA__1_2064 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2064

module FA__1_2067 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2067

module FA__1_2070 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2070

module FA__1_2073 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2073

module FA__1_2076 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2076

module FA__1_2079 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2079

module FA__1_2082 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2082

module HA__1_2085 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2085

module FA__1_2088 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2088

module HA__1_2091 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2091

module FA__1_2094 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2094

module FA__1_2097 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2097

module FA__1_2100 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2100

module HA__1_2103 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2103

module HA__1_2106 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2106

module HA__1_2109 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2109

module HA__1_2112 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2112

module HA__1_2115 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2115

module HA__1_2118 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2118

module HA__1_2121 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2121

module FA__1_2124 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2124

module FA__1_2127 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2127

module FA__1_2130 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2130

module FA__1_2133 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2133

module HA__1_2136 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_2136

module FA__1_2139 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2139

module FA__1_2142 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2142

module FA__1_2145 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2145

module FA__1_2148 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2148

module FA__1_2151 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2151

module WTM8__1_2152 (A_7_PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_7_PP_0;
wire spw_n27;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (spw_n27), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (spw_n27), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (spw_n27), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (spw_n27), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_1965 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_1968 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_1971 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_1974 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_1977 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_1980 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_1983 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_1986 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_1989 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_1992 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_1995 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_1998 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_2001 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_2004 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_2007 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_2010 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_2013 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_2016 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_2019 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_2022 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_2025 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_2028 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_2031 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_2034 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_2037 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_2040 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_2043 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_2046 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_2049 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_2052 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_2055 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_2058 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_2061 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_2064 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_2067 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_2070 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_2073 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_2076 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_2079 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_2082 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_2085 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_2088 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_2091 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_2094 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_2097 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_2100 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_2103 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_2106 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_2109 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_2112 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_2115 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_2118 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_2121 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_2124 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_2127 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_2130 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_2133 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_2136 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_2139 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_2142 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_2145 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_2148 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_2151 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));
BUF_X1 spw__L4_c4_c1 (.Z (spw_n27), .A (A_7_PP_0));

endmodule //WTM8__1_2152

module FA__1_1711 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_1711

module HA__1_1714 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1714

module FA__1_1717 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1717

module FA__1_1720 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1720

module HA__1_1723 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1723

module FA__1_1726 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1726

module FA__1_1729 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1729

module HA__1_1732 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1732

module FA__1_1735 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1735

module FA__1_1738 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1738

module FA__1_1741 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1741

module HA__1_1744 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1744

module FA__1_1747 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1747

module HA__1_1750 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1750

module FA__1_1753 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1753

module FA__1_1756 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1756

module FA__1_1759 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1759

module FA__1_1762 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1762

module FA__1_1765 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1765

module FA__1_1768 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1768

module FA__1_1771 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1771

module FA__1_1774 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1774

module FA__1_1777 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1777

module FA__1_1780 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1780

module FA__1_1783 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1783

module FA__1_1786 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1786

module FA__1_1789 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1789

module FA__1_1792 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1792

module FA__1_1795 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1795

module FA__1_1798 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1798

module FA__1_1801 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1801

module HA__1_1804 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1804

module FA__1_1807 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1807

module FA__1_1810 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1810

module FA__1_1813 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1813

module FA__1_1816 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1816

module FA__1_1819 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1819

module FA__1_1822 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1822

module FA__1_1825 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1825

module FA__1_1828 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1828

module HA__1_1831 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1831

module FA__1_1834 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1834

module HA__1_1837 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1837

module FA__1_1840 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1840

module FA__1_1843 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1843

module FA__1_1846 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1846

module HA__1_1849 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1849

module HA__1_1852 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1852

module HA__1_1855 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1855

module HA__1_1858 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1858

module HA__1_1861 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1861

module HA__1_1864 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1864

module HA__1_1867 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1867

module FA__1_1870 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1870

module FA__1_1873 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1873

module FA__1_1876 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1876

module FA__1_1879 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1879

module HA__1_1882 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1882

module FA__1_1885 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1885

module FA__1_1888 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1888

module FA__1_1891 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1891

module FA__1_1894 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1894

module FA__1_1897 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1897

module WTM8__1_1898 (A_5_PP_0, A_6_PP_0, A_7_PP_0, A_7_PP_1, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_5_PP_0;
input A_6_PP_0;
input A_7_PP_0;
input A_7_PP_1;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A_7_PP_1), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A_6_PP_0), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A_5_PP_0), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A_7_PP_1), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A_6_PP_0), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A_5_PP_0), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A_7_PP_1), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A_6_PP_0), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A_5_PP_0), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A_7_PP_0), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A_5_PP_0), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A_7_PP_0), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A_5_PP_0), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A_7_PP_0), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A_5_PP_0), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_1711 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_1714 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_1717 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_1720 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_1723 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_1726 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_1729 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_1732 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_1735 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_1738 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_1741 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_1744 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_1747 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_1750 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_1753 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_1756 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_1759 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_1762 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_1765 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_1768 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_1771 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_1774 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_1777 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_1780 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_1783 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_1786 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_1789 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_1792 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_1795 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_1798 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_1801 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_1804 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_1807 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_1810 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_1813 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_1816 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_1819 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_1822 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_1825 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_1828 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_1831 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_1834 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_1837 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_1840 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_1843 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_1846 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_1849 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_1852 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_1855 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_1858 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_1861 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_1864 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_1867 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_1870 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_1873 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_1876 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_1879 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_1882 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_1885 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_1888 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_1891 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_1894 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_1897 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__1_1898

module FA__1_3084 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3084

module FA__1_3087 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3087

module FA__1_3090 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3090

module FA__1_3093 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3093

module FA__1_3096 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3096

module FA__1_3099 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3099

module FA__1_3102 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3102

module FA__1_3105 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_3105

module FA__1_3108 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3108

module FA__1_3111 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3111

module FA__1_3114 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3114

module FA__1_3117 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3117

module FA__1_3120 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3120

module FA__1_3123 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3123

module FA__1_3126 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_3126

module FA__1_3129 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_3129

module adder64__1_3178 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;
wire \carry[23] ;
wire \carry[22] ;
wire \carry[21] ;
wire \carry[20] ;
wire \carry[19] ;
wire \carry[18] ;
wire \carry[17] ;
wire \carry[16] ;


FA__1_3084 genblk1_31_F (.carry (z[32]), .sum (z[31]), .b (y[31]), .cin (\carry[30] ));
FA__1_3087 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .b (y[30]), .cin (\carry[29] ));
FA__1_3090 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .b (y[29]), .cin (\carry[28] ));
FA__1_3093 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .b (y[28]), .cin (\carry[27] ));
FA__1_3096 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .b (y[27]), .cin (\carry[26] ));
FA__1_3099 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .b (y[26]), .cin (\carry[25] ));
FA__1_3102 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .b (y[25]), .cin (\carry[24] ));
FA__1_3105 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .b (y[24]), .cin (\carry[23] ));
FA__1_3108 genblk1_23_F (.carry (\carry[23] ), .sum (z[23]), .a (x[23]), .b (y[23]), .cin (\carry[22] ));
FA__1_3111 genblk1_22_F (.carry (\carry[22] ), .sum (z[22]), .a (x[22]), .b (y[22]), .cin (\carry[21] ));
FA__1_3114 genblk1_21_F (.carry (\carry[21] ), .sum (z[21]), .a (x[21]), .b (y[21]), .cin (\carry[20] ));
FA__1_3117 genblk1_20_F (.carry (\carry[20] ), .sum (z[20]), .a (x[20]), .b (y[20]), .cin (\carry[19] ));
FA__1_3120 genblk1_19_F (.carry (\carry[19] ), .sum (z[19]), .a (x[19]), .b (y[19]), .cin (\carry[18] ));
FA__1_3123 genblk1_18_F (.carry (\carry[18] ), .sum (z[18]), .a (x[18]), .b (y[18]), .cin (\carry[17] ));
FA__1_3126 genblk1_17_F (.carry (\carry[17] ), .sum (z[17]), .a (x[17]), .b (y[17]), .cin (\carry[16] ));
FA__1_3129 genblk1_16_F (.carry (\carry[16] ), .sum (z[16]), .a (x[16]), .b (y[16]));

endmodule //adder64__1_3178

module FA__1_1457 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_1457

module HA__1_1460 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1460

module FA__1_1463 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1463

module FA__1_1466 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1466

module HA__1_1469 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1469

module FA__1_1472 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1472

module FA__1_1475 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1475

module HA__1_1478 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1478

module FA__1_1481 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1481

module FA__1_1484 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1484

module FA__1_1487 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1487

module HA__1_1490 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1490

module FA__1_1493 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1493

module HA__1_1496 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1496

module FA__1_1499 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1499

module FA__1_1502 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1502

module FA__1_1505 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1505

module FA__1_1508 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1508

module FA__1_1511 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1511

module FA__1_1514 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1514

module FA__1_1517 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1517

module FA__1_1520 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1520

module FA__1_1523 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1523

module FA__1_1526 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1526

module FA__1_1529 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1529

module FA__1_1532 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1532

module FA__1_1535 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1535

module FA__1_1538 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1538

module FA__1_1541 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1541

module FA__1_1544 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1544

module FA__1_1547 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1547

module HA__1_1550 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1550

module FA__1_1553 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1553

module FA__1_1556 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1556

module FA__1_1559 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1559

module FA__1_1562 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1562

module FA__1_1565 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1565

module FA__1_1568 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1568

module FA__1_1571 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1571

module FA__1_1574 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1574

module HA__1_1577 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1577

module FA__1_1580 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1580

module HA__1_1583 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1583

module FA__1_1586 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1586

module FA__1_1589 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1589

module FA__1_1592 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1592

module HA__1_1595 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1595

module HA__1_1598 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1598

module HA__1_1601 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1601

module HA__1_1604 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1604

module HA__1_1607 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1607

module HA__1_1610 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1610

module HA__1_1613 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1613

module FA__1_1616 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1616

module FA__1_1619 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1619

module FA__1_1622 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1622

module FA__1_1625 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1625

module HA__1_1628 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1628

module FA__1_1631 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1631

module FA__1_1634 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1634

module FA__1_1637 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1637

module FA__1_1640 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1640

module FA__1_1643 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1643

module WTM8__1_1644 (B_7_PP_0, B_5_PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input B_7_PP_0;
input B_5_PP_0;
wire spw_n22;
wire spw_n50;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (spw_n50));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (spw_n50));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (spw_n50));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (spw_n22));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (spw_n22));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (spw_n22));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_1457 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_1460 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_1463 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_1466 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_1469 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_1472 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_1475 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_1478 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_1481 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_1484 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_1487 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_1490 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_1493 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_1496 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_1499 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_1502 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_1505 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_1508 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_1511 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_1514 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_1517 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_1520 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_1523 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_1526 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_1529 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_1532 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_1535 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_1538 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_1541 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_1544 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_1547 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_1550 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_1553 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_1556 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_1559 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_1562 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_1565 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_1568 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_1571 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_1574 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_1577 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_1580 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_1583 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_1586 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_1589 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_1592 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_1595 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_1598 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_1601 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_1604 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_1607 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_1610 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_1613 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_1616 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_1619 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_1622 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_1625 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_1628 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_1631 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_1634 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_1637 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_1640 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_1643 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));
BUF_X1 spw__L4_c4_c1 (.Z (spw_n22), .A (B_7_PP_0));
BUF_X1 spw__L5_c8_c4 (.Z (spw_n50), .A (B_5_PP_0));

endmodule //WTM8__1_1644

module FA__1_1203 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_1203

module HA__1_1206 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1206

module FA__1_1209 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1209

module FA__1_1212 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1212

module HA__1_1215 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1215

module FA__1_1218 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1218

module FA__1_1221 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1221

module HA__1_1224 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1224

module FA__1_1227 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1227

module FA__1_1230 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1230

module FA__1_1233 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1233

module HA__1_1236 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1236

module FA__1_1239 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1239

module HA__1_1242 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1242

module FA__1_1245 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1245

module FA__1_1248 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1248

module FA__1_1251 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1251

module FA__1_1254 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1254

module FA__1_1257 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1257

module FA__1_1260 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1260

module FA__1_1263 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1263

module FA__1_1266 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1266

module FA__1_1269 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1269

module FA__1_1272 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1272

module FA__1_1275 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1275

module FA__1_1278 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1278

module FA__1_1281 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1281

module FA__1_1284 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1284

module FA__1_1287 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1287

module FA__1_1290 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1290

module FA__1_1293 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1293

module HA__1_1296 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1296

module FA__1_1299 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1299

module FA__1_1302 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1302

module FA__1_1305 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1305

module FA__1_1308 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1308

module FA__1_1311 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1311

module FA__1_1314 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1314

module FA__1_1317 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1317

module FA__1_1320 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1320

module HA__1_1323 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1323

module FA__1_1326 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1326

module HA__1_1329 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1329

module FA__1_1332 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1332

module FA__1_1335 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1335

module FA__1_1338 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1338

module HA__1_1341 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1341

module HA__1_1344 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1344

module HA__1_1347 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1347

module HA__1_1350 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1350

module HA__1_1353 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1353

module HA__1_1356 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1356

module HA__1_1359 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1359

module FA__1_1362 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1362

module FA__1_1365 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1365

module FA__1_1368 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1368

module FA__1_1371 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1371

module HA__1_1374 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1374

module FA__1_1377 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1377

module FA__1_1380 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1380

module FA__1_1383 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1383

module FA__1_1386 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1386

module FA__1_1389 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1389

module WTM8__1_1390 (A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_1203 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_1206 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_1209 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_1212 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_1215 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_1218 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_1221 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_1224 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_1227 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_1230 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_1233 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_1236 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_1239 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_1242 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_1245 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_1248 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_1251 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_1254 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_1257 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_1260 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_1263 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_1266 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_1269 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_1272 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_1275 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_1278 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_1281 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_1284 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_1287 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_1290 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_1293 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_1296 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_1299 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_1302 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_1305 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_1308 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_1311 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_1314 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_1317 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_1320 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_1323 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_1326 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_1329 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_1332 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_1335 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_1338 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_1341 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_1344 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_1347 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_1350 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_1353 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_1356 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_1359 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_1362 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_1365 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_1368 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_1371 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_1374 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_1377 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_1380 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_1383 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_1386 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_1389 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__1_1390

module FA__1_2864 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2864

module FA__1_2867 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2867

module FA__1_2870 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2870

module FA__1_2873 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2873

module FA__1_2876 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2876

module FA__1_2879 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2879

module FA__1_2882 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2882

module FA__1_2885 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2885

module FA__1_2888 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2888

module FA__1_2891 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2891

module FA__1_2894 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2894

module FA__1_2897 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2897

module FA__1_2900 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2900

module FA__1_2903 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2903

module FA__1_2906 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2906

module FA__1_2909 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2909

module FA__1_2912 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2912

module FA__1_2915 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2915

module FA__1_2918 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2918

module FA__1_2921 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2921

module FA__1_2924 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2924

module FA__1_2927 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2927

module FA__1_2930 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2930

module FA__1_2933 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2933

module FA__1_2936 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X2 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_2936

module adder64__1_2985 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;
wire \carry[23] ;
wire \carry[22] ;
wire \carry[21] ;
wire \carry[20] ;
wire \carry[19] ;
wire \carry[18] ;
wire \carry[17] ;
wire \carry[16] ;


FA__1_2864 genblk1_40_F (.carry (z[41]), .sum (z[40]), .b (y[40]), .cin (\carry[39] ));
FA__1_2867 genblk1_39_F (.carry (\carry[39] ), .sum (z[39]), .b (y[39]), .cin (\carry[38] ));
FA__1_2870 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .b (y[38]), .cin (\carry[37] ));
FA__1_2873 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .b (y[37]), .cin (\carry[36] ));
FA__1_2876 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .b (y[36]), .cin (\carry[35] ));
FA__1_2879 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .b (y[35]), .cin (\carry[34] ));
FA__1_2882 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .b (y[34]), .cin (\carry[33] ));
FA__1_2885 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .b (y[33]), .cin (\carry[32] ));
FA__1_2888 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .b (y[32]), .cin (\carry[31] ));
FA__1_2891 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .b (y[31]), .cin (\carry[30] ));
FA__1_2894 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .b (y[30]), .cin (\carry[29] ));
FA__1_2897 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .b (y[29]), .cin (\carry[28] ));
FA__1_2900 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .b (y[28]), .cin (\carry[27] ));
FA__1_2903 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .b (y[27]), .cin (\carry[26] ));
FA__1_2906 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .b (y[26]), .cin (\carry[25] ));
FA__1_2909 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .b (y[25]), .cin (\carry[24] ));
FA__1_2912 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24])
    , .cin (\carry[23] ));
FA__1_2915 genblk1_23_F (.carry (\carry[23] ), .sum (z[23]), .a (x[23]), .b (y[23])
    , .cin (\carry[22] ));
FA__1_2918 genblk1_22_F (.carry (\carry[22] ), .sum (z[22]), .a (x[22]), .b (y[22])
    , .cin (\carry[21] ));
FA__1_2921 genblk1_21_F (.carry (\carry[21] ), .sum (z[21]), .a (x[21]), .b (y[21])
    , .cin (\carry[20] ));
FA__1_2924 genblk1_20_F (.carry (\carry[20] ), .sum (z[20]), .a (x[20]), .b (y[20])
    , .cin (\carry[19] ));
FA__1_2927 genblk1_19_F (.carry (\carry[19] ), .sum (z[19]), .a (x[19]), .b (y[19])
    , .cin (\carry[18] ));
FA__1_2930 genblk1_18_F (.carry (\carry[18] ), .sum (z[18]), .a (x[18]), .b (y[18])
    , .cin (\carry[17] ));
FA__1_2933 genblk1_17_F (.carry (\carry[17] ), .sum (z[17]), .a (x[17]), .b (y[17])
    , .cin (\carry[16] ));
FA__1_2936 genblk1_16_F (.carry (\carry[16] ), .sum (z[16]), .a (x[16]), .b (y[16]));

endmodule //adder64__1_2985

module FA__1_2674 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2674

module FA__1_2677 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2677

module FA__1_2680 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2680

module FA__1_2683 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2683

module FA__1_2686 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2686

module FA__1_2689 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2689

module FA__1_2692 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2692

module FA__1_2695 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2695

module FA__1_2698 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2698

module FA__1_2701 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2701

module FA__1_2704 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2704

module FA__1_2707 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2707

module FA__1_2710 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2710

module FA__1_2713 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2713

module FA__1_2716 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2716

module FA__1_2719 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_2719

module adder64__1_2792 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;


FA__1_2674 genblk1_39_F (.carry (z[40]), .sum (z[39]), .b (y[39]), .cin (\carry[38] ));
FA__1_2677 genblk1_38_F (.carry (\carry[38] ), .sum (z[38]), .b (y[38]), .cin (\carry[37] ));
FA__1_2680 genblk1_37_F (.carry (\carry[37] ), .sum (z[37]), .b (y[37]), .cin (\carry[36] ));
FA__1_2683 genblk1_36_F (.carry (\carry[36] ), .sum (z[36]), .b (y[36]), .cin (\carry[35] ));
FA__1_2686 genblk1_35_F (.carry (\carry[35] ), .sum (z[35]), .b (y[35]), .cin (\carry[34] ));
FA__1_2689 genblk1_34_F (.carry (\carry[34] ), .sum (z[34]), .b (y[34]), .cin (\carry[33] ));
FA__1_2692 genblk1_33_F (.carry (\carry[33] ), .sum (z[33]), .b (y[33]), .cin (\carry[32] ));
FA__1_2695 genblk1_32_F (.carry (\carry[32] ), .sum (z[32]), .b (y[32]), .cin (\carry[31] ));
FA__1_2698 genblk1_31_F (.carry (\carry[31] ), .sum (z[31]), .a (x[31]), .b (y[31]), .cin (\carry[30] ));
FA__1_2701 genblk1_30_F (.carry (\carry[30] ), .sum (z[30]), .a (x[30]), .b (y[30]), .cin (\carry[29] ));
FA__1_2704 genblk1_29_F (.carry (\carry[29] ), .sum (z[29]), .a (x[29]), .b (y[29]), .cin (\carry[28] ));
FA__1_2707 genblk1_28_F (.carry (\carry[28] ), .sum (z[28]), .a (x[28]), .b (y[28]), .cin (\carry[27] ));
FA__1_2710 genblk1_27_F (.carry (\carry[27] ), .sum (z[27]), .a (x[27]), .b (y[27]), .cin (\carry[26] ));
FA__1_2713 genblk1_26_F (.carry (\carry[26] ), .sum (z[26]), .a (x[26]), .b (y[26]), .cin (\carry[25] ));
FA__1_2716 genblk1_25_F (.carry (\carry[25] ), .sum (z[25]), .a (x[25]), .b (y[25]), .cin (\carry[24] ));
FA__1_2719 genblk1_24_F (.carry (\carry[24] ), .sum (z[24]), .a (x[24]), .b (y[24]));

endmodule //adder64__1_2792

module FA__1_949 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_949

module HA__1_952 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_952

module FA__1_955 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_955

module FA__1_958 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_958

module HA__1_961 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_961

module FA__1_964 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_964

module FA__1_967 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_967

module HA__1_970 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_970

module FA__1_973 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_973

module FA__1_976 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_976

module FA__1_979 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_979

module HA__1_982 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_982

module FA__1_985 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_985

module HA__1_988 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_988

module FA__1_991 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_991

module FA__1_994 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_994

module FA__1_997 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_997

module FA__1_1000 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1000

module FA__1_1003 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1003

module FA__1_1006 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1006

module FA__1_1009 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1009

module FA__1_1012 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1012

module FA__1_1015 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1015

module FA__1_1018 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1018

module FA__1_1021 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1021

module FA__1_1024 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1024

module FA__1_1027 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1027

module FA__1_1030 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1030

module FA__1_1033 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1033

module FA__1_1036 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1036

module FA__1_1039 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1039

module HA__1_1042 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1042

module FA__1_1045 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1045

module FA__1_1048 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1048

module FA__1_1051 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1051

module FA__1_1054 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1054

module FA__1_1057 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1057

module FA__1_1060 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1060

module FA__1_1063 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1063

module FA__1_1066 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1066

module HA__1_1069 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1069

module FA__1_1072 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1072

module HA__1_1075 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1075

module FA__1_1078 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1078

module FA__1_1081 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1081

module FA__1_1084 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1084

module HA__1_1087 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1087

module HA__1_1090 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1090

module HA__1_1093 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1093

module HA__1_1096 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1096

module HA__1_1099 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1099

module HA__1_1102 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1102

module HA__1_1105 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1105

module FA__1_1108 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1108

module FA__1_1111 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1111

module FA__1_1114 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1114

module FA__1_1117 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1117

module HA__1_1120 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_1120

module FA__1_1123 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1123

module FA__1_1126 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1126

module FA__1_1129 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1129

module FA__1_1132 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1132

module FA__1_1135 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_1135

module WTM8__1_1136 (A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_949 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_952 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_955 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_958 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_961 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_964 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_967 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_970 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_973 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_976 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_979 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_982 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_985 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_988 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_991 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_994 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_997 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_1000 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_1003 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_1006 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_1009 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_1012 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_1015 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_1018 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_1021 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_1024 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_1027 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_1030 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_1033 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_1036 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_1039 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_1042 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_1045 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_1048 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_1051 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_1054 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_1057 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_1060 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_1063 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_1066 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_1069 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_1072 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_1075 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_1078 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_1081 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_1084 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_1087 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_1090 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_1093 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_1096 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_1099 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_1102 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_1105 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_1108 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_1111 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_1114 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_1117 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_1120 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_1123 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_1126 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_1129 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_1132 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_1135 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__1_1136

module FA__1_695 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_695

module HA__1_698 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_698

module FA__1_701 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_701

module FA__1_704 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_704

module HA__1_707 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_707

module FA__1_710 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_710

module FA__1_713 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_713

module HA__1_716 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_716

module FA__1_719 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_719

module FA__1_722 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_722

module FA__1_725 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_725

module HA__1_728 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_728

module FA__1_731 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_731

module HA__1_734 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_734

module FA__1_737 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_737

module FA__1_740 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_740

module FA__1_743 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_743

module FA__1_746 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_746

module FA__1_749 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_749

module FA__1_752 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_752

module FA__1_755 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_755

module FA__1_758 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_758

module FA__1_761 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_761

module FA__1_764 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_764

module FA__1_767 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_767

module FA__1_770 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_770

module FA__1_773 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_773

module FA__1_776 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_776

module FA__1_779 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_779

module FA__1_782 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_782

module FA__1_785 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_785

module HA__1_788 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_788

module FA__1_791 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_791

module FA__1_794 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_794

module FA__1_797 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_797

module FA__1_800 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_800

module FA__1_803 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_803

module FA__1_806 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_806

module FA__1_809 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_809

module FA__1_812 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_812

module HA__1_815 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_815

module FA__1_818 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_818

module HA__1_821 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_821

module FA__1_824 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_824

module FA__1_827 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_827

module FA__1_830 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_830

module HA__1_833 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_833

module HA__1_836 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_836

module HA__1_839 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_839

module HA__1_842 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_842

module HA__1_845 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_845

module HA__1_848 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_848

module HA__1_851 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_851

module FA__1_854 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_854

module FA__1_857 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_857

module FA__1_860 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_860

module FA__1_863 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_863

module HA__1_866 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_866

module FA__1_869 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_869

module FA__1_872 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_872

module FA__1_875 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_875

module FA__1_878 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_878

module FA__1_881 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_881

module WTM8__1_882 (A_7_PP_0, A_6_PP_0, A_5_PP_0, A_5_PP_1, A_6_PP_0PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input A_7_PP_0;
input A_6_PP_0;
input A_5_PP_0;
input A_5_PP_1;
input A_6_PP_0PP_0;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X1 i_0_51 (.ZN (n_157), .A1 (A_7_PP_0), .A2 (B[0]));
AND2_X1 i_0_50 (.ZN (n_156), .A1 (A_6_PP_0PP_0), .A2 (B[0]));
AND2_X1 i_0_49 (.ZN (n_155), .A1 (A_5_PP_1), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A_7_PP_0), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A_6_PP_0PP_0), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A_5_PP_0), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A_6_PP_0), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A_5_PP_0), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B[5]));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B[5]));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B[5]));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B[5]));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B[5]));
AND2_X1 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B[5]));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_695 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_698 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_701 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_704 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_707 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_710 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_713 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_716 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_719 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_722 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_725 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_728 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_731 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_734 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_737 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_740 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_743 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_746 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_749 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_752 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_755 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_758 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_761 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_764 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_767 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_770 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_773 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_776 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_779 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_782 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_785 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_788 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_791 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_794 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_797 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_800 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_803 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_806 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_809 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_812 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_815 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_818 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_821 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_824 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_827 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_830 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_833 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_836 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_839 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_842 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_845 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_848 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_851 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_854 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_857 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_860 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_863 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_866 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_869 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_872 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_875 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_878 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_881 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__1_882

module FA__1_2529 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2529

module FA__1_2532 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2532

module FA__1_2535 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2535

module FA__1_2538 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2538

module FA__1_2541 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2541

module FA__1_2544 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2544

module FA__1_2547 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X2 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2547

module FA__1_2550 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X2 i_0_1 (.ZN (carry), .A1 (b), .A2 (cin));
XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (b));

endmodule //FA__1_2550

module FA__1_2553 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2553

module FA__1_2556 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2556

module FA__1_2559 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2559

module FA__1_2562 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X4 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2562

module FA__1_2565 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2565

module FA__1_2568 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2568

module FA__1_2571 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_2571

module FA__1_2574 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;


AND2_X1 i_0_1 (.ZN (carry), .A1 (b), .A2 (a));
XOR2_X1 i_0_0 (.Z (sum), .A (a), .B (b));

endmodule //FA__1_2574

module adder64__1_2599 (x, y, z, C);

output C;
output [63:0] z;
input [63:0] x;
input [63:0] y;
wire \carry[22] ;
wire \carry[21] ;
wire \carry[20] ;
wire \carry[19] ;
wire \carry[18] ;
wire \carry[17] ;
wire \carry[16] ;
wire \carry[15] ;
wire \carry[14] ;
wire \carry[13] ;
wire \carry[12] ;
wire \carry[11] ;
wire \carry[10] ;
wire \carry[9] ;
wire \carry[8] ;


FA__1_2529 genblk1_23_F (.carry (z[24]), .sum (z[23]), .b (y[23]), .cin (\carry[22] ));
FA__1_2532 genblk1_22_F (.carry (\carry[22] ), .sum (z[22]), .b (y[22]), .cin (\carry[21] ));
FA__1_2535 genblk1_21_F (.carry (\carry[21] ), .sum (z[21]), .b (y[21]), .cin (\carry[20] ));
FA__1_2538 genblk1_20_F (.carry (\carry[20] ), .sum (z[20]), .b (y[20]), .cin (\carry[19] ));
FA__1_2541 genblk1_19_F (.carry (\carry[19] ), .sum (z[19]), .b (y[19]), .cin (\carry[18] ));
FA__1_2544 genblk1_18_F (.carry (\carry[18] ), .sum (z[18]), .b (y[18]), .cin (\carry[17] ));
FA__1_2547 genblk1_17_F (.carry (\carry[17] ), .sum (z[17]), .b (y[17]), .cin (\carry[16] ));
FA__1_2550 genblk1_16_F (.carry (\carry[16] ), .sum (z[16]), .b (y[16]), .cin (\carry[15] ));
FA__1_2553 genblk1_15_F (.carry (\carry[15] ), .sum (z[15]), .a (x[15]), .b (y[15])
    , .cin (\carry[14] ));
FA__1_2556 genblk1_14_F (.carry (\carry[14] ), .sum (z[14]), .a (x[14]), .b (y[14])
    , .cin (\carry[13] ));
FA__1_2559 genblk1_13_F (.carry (\carry[13] ), .sum (z[13]), .a (x[13]), .b (y[13])
    , .cin (\carry[12] ));
FA__1_2562 genblk1_12_F (.carry (\carry[12] ), .sum (z[12]), .a (x[12]), .b (y[12])
    , .cin (\carry[11] ));
FA__1_2565 genblk1_11_F (.carry (\carry[11] ), .sum (z[11]), .a (x[11]), .b (y[11])
    , .cin (\carry[10] ));
FA__1_2568 genblk1_10_F (.carry (\carry[10] ), .sum (z[10]), .a (x[10]), .b (y[10]), .cin (\carry[9] ));
FA__1_2571 genblk1_9_F (.carry (\carry[9] ), .sum (z[9]), .a (x[9]), .b (y[9]), .cin (\carry[8] ));
FA__1_2574 genblk1_8_F (.carry (\carry[8] ), .sum (z[8]), .a (x[8]), .b (y[8]));

endmodule //adder64__1_2599

module FA__1_441 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;


XNOR2_X2 i_0_1 (.ZN (sum), .A (n_0_0), .B (b));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (a), .B (cin));

endmodule //FA__1_441

module HA__1_444 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_444

module FA__1_447 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_447

module FA__1_450 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_450

module HA__1_453 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_453

module FA__1_456 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_456

module FA__1_459 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_459

module HA__1_462 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_462

module FA__1_465 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_465

module FA__1_468 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_468

module FA__1_471 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_471

module HA__1_474 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_474

module FA__1_477 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_477

module HA__1_480 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_480

module FA__1_483 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_483

module FA__1_486 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_486

module FA__1_489 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_489

module FA__1_492 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_492

module FA__1_495 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_495

module FA__1_498 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_498

module FA__1_501 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_501

module FA__1_504 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_504

module FA__1_507 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_507

module FA__1_510 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_510

module FA__1_513 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_513

module FA__1_516 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_516

module FA__1_519 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_519

module FA__1_522 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_522

module FA__1_525 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_525

module FA__1_528 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_528

module FA__1_531 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_531

module HA__1_534 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_534

module FA__1_537 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_537

module FA__1_540 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_540

module FA__1_543 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_543

module FA__1_546 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_546

module FA__1_549 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_549

module FA__1_552 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_552

module FA__1_555 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_555

module FA__1_558 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X2 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_558

module HA__1_561 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X2 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_561

module FA__1_564 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_564

module HA__1_567 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_567

module FA__1_570 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_570

module FA__1_573 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_573

module FA__1_576 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_576

module HA__1_579 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X2 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_579

module HA__1_582 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_582

module HA__1_585 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_585

module HA__1_588 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_588

module HA__1_591 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_591

module HA__1_594 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_594

module HA__1_597 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_597

module FA__1_600 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_600

module FA__1_603 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_603

module FA__1_606 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_606

module FA__1_609 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_609

module HA__1_612 (a, b, s, c);

output c;
output s;
input a;
input b;


AND2_X1 i_0_1 (.ZN (c), .A1 (a), .A2 (b));
XOR2_X1 i_0_0 (.Z (s), .A (a), .B (b));

endmodule //HA__1_612

module FA__1_615 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_615

module FA__1_618 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_618

module FA__1_621 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_621

module FA__1_624 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X1 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_624

module FA__1_627 (a, b, cin, sum, carry);

output carry;
output sum;
input a;
input b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (a));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (cin), .B (a));
XNOR2_X2 i_0_2 (.ZN (sum), .A (b), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (b), .B1 (cin), .B2 (a));
NAND2_X1 i_0_0 (.ZN (carry), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__1_627

module WTM8__1_628 (B_5_PP_0, A, B, Result);

output [15:0] Result;
input [7:0] A;
input [7:0] B;
input B_5_PP_0;
wire C;
wire S;
wire P;
wire n_155;
wire n_147;
wire n_139;
wire n_161;
wire n_154;
wire n_146;
wire n_1;
wire n_0;
wire n_131;
wire n_123;
wire n_116;
wire n_3;
wire n_2;
wire n_5;
wire n_4;
wire n_160;
wire n_153;
wire n_145;
wire n_7;
wire n_6;
wire n_138;
wire n_130;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_13;
wire n_12;
wire n_159;
wire n_152;
wire n_144;
wire n_15;
wire n_14;
wire n_137;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_21;
wire n_20;
wire n_158;
wire n_151;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_156;
wire n_148;
wire n_140;
wire n_28;
wire n_27;
wire n_132;
wire n_124;
wire n_117;
wire n_30;
wire n_29;
wire n_32;
wire n_31;
wire n_162;
wire n_34;
wire n_33;
wire n_36;
wire n_35;
wire n_38;
wire n_37;
wire n_39;
wire n_157;
wire n_149;
wire n_141;
wire n_41;
wire n_40;
wire n_133;
wire n_125;
wire n_118;
wire n_43;
wire n_42;
wire n_45;
wire n_44;
wire n_163;
wire n_108;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_52;
wire n_150;
wire n_142;
wire n_54;
wire n_53;
wire n_134;
wire n_126;
wire n_120;
wire n_56;
wire n_55;
wire n_58;
wire n_57;
wire n_164;
wire n_109;
wire n_60;
wire n_59;
wire n_62;
wire n_61;
wire n_64;
wire n_63;
wire n_65;
wire n_143;
wire n_135;
wire n_127;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_119;
wire n_165;
wire n_110;
wire n_71;
wire n_70;
wire n_73;
wire n_72;
wire n_75;
wire n_74;
wire n_76;
wire n_136;
wire n_128;
wire n_121;
wire n_78;
wire n_77;
wire n_166;
wire n_111;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_83;
wire n_85;
wire n_129;
wire n_87;
wire n_86;
wire n_167;
wire n_112;
wire n_89;
wire n_88;
wire n_91;
wire n_90;
wire n_93;
wire n_92;
wire n_94;
wire n_122;
wire n_168;
wire n_113;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_100;
wire n_99;
wire n_101;
wire n_169;
wire n_114;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_106;
wire n_115;
wire n_107;


AND2_X1 i_0_63 (.ZN (n_169), .A1 (A[7]), .A2 (B[6]));
AND2_X1 i_0_62 (.ZN (n_168), .A1 (A[6]), .A2 (B[6]));
AND2_X1 i_0_61 (.ZN (n_167), .A1 (A[5]), .A2 (B[6]));
AND2_X1 i_0_60 (.ZN (n_166), .A1 (A[4]), .A2 (B[6]));
AND2_X1 i_0_59 (.ZN (n_165), .A1 (A[3]), .A2 (B[6]));
AND2_X1 i_0_58 (.ZN (n_164), .A1 (A[2]), .A2 (B[6]));
AND2_X1 i_0_57 (.ZN (n_163), .A1 (A[1]), .A2 (B[6]));
AND2_X1 i_0_56 (.ZN (n_162), .A1 (A[0]), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_161), .A1 (A[4]), .A2 (B[0]));
AND2_X1 i_0_54 (.ZN (n_160), .A1 (A[3]), .A2 (B[0]));
AND2_X1 i_0_53 (.ZN (n_159), .A1 (A[2]), .A2 (B[0]));
AND2_X1 i_0_52 (.ZN (n_158), .A1 (A[1]), .A2 (B[0]));
AND2_X4 i_0_51 (.ZN (n_157), .A1 (A[7]), .A2 (B[0]));
AND2_X4 i_0_50 (.ZN (n_156), .A1 (A[6]), .A2 (B[0]));
AND2_X4 i_0_49 (.ZN (n_155), .A1 (A[5]), .A2 (B[0]));
AND2_X1 i_0_48 (.ZN (n_154), .A1 (A[3]), .A2 (B[1]));
AND2_X1 i_0_47 (.ZN (n_153), .A1 (A[2]), .A2 (B[1]));
AND2_X1 i_0_46 (.ZN (n_152), .A1 (A[1]), .A2 (B[1]));
AND2_X1 i_0_45 (.ZN (n_151), .A1 (A[0]), .A2 (B[1]));
AND2_X1 i_0_44 (.ZN (n_150), .A1 (A[7]), .A2 (B[1]));
AND2_X1 i_0_43 (.ZN (n_149), .A1 (A[6]), .A2 (B[1]));
AND2_X1 i_0_42 (.ZN (n_148), .A1 (A[5]), .A2 (B[1]));
AND2_X1 i_0_41 (.ZN (n_147), .A1 (A[4]), .A2 (B[1]));
AND2_X1 i_0_40 (.ZN (n_146), .A1 (A[2]), .A2 (B[2]));
AND2_X1 i_0_39 (.ZN (n_145), .A1 (A[1]), .A2 (B[2]));
AND2_X1 i_0_38 (.ZN (n_144), .A1 (A[0]), .A2 (B[2]));
AND2_X1 i_0_37 (.ZN (n_143), .A1 (A[7]), .A2 (B[2]));
AND2_X1 i_0_36 (.ZN (n_142), .A1 (A[6]), .A2 (B[2]));
AND2_X1 i_0_35 (.ZN (n_141), .A1 (A[5]), .A2 (B[2]));
AND2_X1 i_0_34 (.ZN (n_140), .A1 (A[4]), .A2 (B[2]));
AND2_X1 i_0_33 (.ZN (n_139), .A1 (A[3]), .A2 (B[2]));
AND2_X1 i_0_32 (.ZN (n_138), .A1 (A[1]), .A2 (B[3]));
AND2_X1 i_0_31 (.ZN (n_137), .A1 (A[0]), .A2 (B[3]));
AND2_X1 i_0_30 (.ZN (n_136), .A1 (A[7]), .A2 (B[3]));
AND2_X1 i_0_29 (.ZN (n_135), .A1 (A[6]), .A2 (B[3]));
AND2_X1 i_0_28 (.ZN (n_134), .A1 (A[5]), .A2 (B[3]));
AND2_X1 i_0_27 (.ZN (n_133), .A1 (A[4]), .A2 (B[3]));
AND2_X1 i_0_26 (.ZN (n_132), .A1 (A[3]), .A2 (B[3]));
AND2_X1 i_0_25 (.ZN (n_131), .A1 (A[2]), .A2 (B[3]));
AND2_X1 i_0_24 (.ZN (n_130), .A1 (A[0]), .A2 (B[4]));
AND2_X1 i_0_23 (.ZN (n_129), .A1 (A[7]), .A2 (B[4]));
AND2_X1 i_0_22 (.ZN (n_128), .A1 (A[6]), .A2 (B[4]));
AND2_X1 i_0_21 (.ZN (n_127), .A1 (A[5]), .A2 (B[4]));
AND2_X1 i_0_20 (.ZN (n_126), .A1 (A[4]), .A2 (B[4]));
AND2_X1 i_0_19 (.ZN (n_125), .A1 (A[3]), .A2 (B[4]));
AND2_X1 i_0_18 (.ZN (n_124), .A1 (A[2]), .A2 (B[4]));
AND2_X1 i_0_17 (.ZN (n_123), .A1 (A[1]), .A2 (B[4]));
AND2_X1 i_0_16 (.ZN (P), .A1 (A[6]), .A2 (B[5]));
AND2_X1 i_0_15 (.ZN (n_122), .A1 (A[7]), .A2 (B[5]));
AND2_X1 i_0_14 (.ZN (n_121), .A1 (A[5]), .A2 (B_5_PP_0));
AND2_X1 i_0_13 (.ZN (n_120), .A1 (A[3]), .A2 (B_5_PP_0));
AND2_X1 i_0_12 (.ZN (n_119), .A1 (A[4]), .A2 (B_5_PP_0));
AND2_X1 i_0_11 (.ZN (n_118), .A1 (A[2]), .A2 (B_5_PP_0));
AND2_X1 i_0_10 (.ZN (n_117), .A1 (A[1]), .A2 (B_5_PP_0));
AND2_X4 i_0_9 (.ZN (n_116), .A1 (A[0]), .A2 (B_5_PP_0));
AND2_X1 i_0_8 (.ZN (n_115), .A1 (A[7]), .A2 (B[7]));
AND2_X1 i_0_7 (.ZN (n_114), .A1 (A[6]), .A2 (B[7]));
AND2_X1 i_0_6 (.ZN (n_113), .A1 (A[5]), .A2 (B[7]));
AND2_X1 i_0_5 (.ZN (n_112), .A1 (A[4]), .A2 (B[7]));
AND2_X1 i_0_4 (.ZN (n_111), .A1 (A[3]), .A2 (B[7]));
AND2_X1 i_0_3 (.ZN (n_110), .A1 (A[2]), .A2 (B[7]));
AND2_X1 i_0_2 (.ZN (n_109), .A1 (A[1]), .A2 (B[7]));
AND2_X1 i_0_1 (.ZN (n_108), .A1 (A[0]), .A2 (B[7]));
AND2_X1 i_0_0 (.ZN (Result[0]), .A1 (A[0]), .A2 (B[0]));
FA__1_441 F46 (.sum (Result[14]), .a (n_107), .b (n_104), .cin (n_106));
HA__1_444 H14 (.c (Result[15]), .s (n_107), .a (n_115), .b (n_102));
FA__1_447 F45 (.carry (n_106), .sum (Result[13]), .a (n_105), .b (n_99), .cin (n_101));
FA__1_450 F37 (.carry (n_104), .sum (n_105), .a (n_97), .b (n_103), .cin (n_95));
HA__1_453 H5 (.c (n_102), .s (n_103), .a (n_169), .b (n_114));
FA__1_456 F44 (.carry (n_101), .sum (Result[12]), .a (n_100), .b (n_92), .cin (n_94));
FA__1_459 F36 (.carry (n_99), .sum (n_100), .a (n_98), .b (n_88), .cin (n_90));
HA__1_462 H10 (.c (n_97), .s (n_98), .a (n_86), .b (n_96));
FA__1_465 F21 (.carry (n_95), .sum (n_96), .a (n_122), .b (n_168), .cin (n_113));
FA__1_468 F43 (.carry (n_94), .sum (Result[11]), .a (n_93), .b (n_83), .cin (n_85));
FA__1_471 F35 (.carry (n_92), .sum (n_93), .a (n_91), .b (n_81), .cin (n_79));
HA__1_474 H9 (.c (n_90), .s (n_91), .a (n_87), .b (n_89));
FA__1_477 F20 (.carry (n_88), .sum (n_89), .a (n_77), .b (n_167), .cin (n_112));
HA__1_480 H3 (.c (n_86), .s (n_87), .a (n_129), .b (P));
FA__1_483 F42 (.carry (n_85), .sum (Result[10]), .a (n_84), .b (n_74), .cin (n_76));
FA__1_486 F34 (.carry (n_83), .sum (n_84), .a (n_82), .b (n_72), .cin (n_70));
FA__1_489 F30 (.carry (n_81), .sum (n_82), .a (n_78), .b (n_68), .cin (n_80));
FA__1_492 F19 (.carry (n_79), .sum (n_80), .a (n_66), .b (n_166), .cin (n_111));
FA__1_495 F11 (.carry (n_77), .sum (n_78), .a (n_136), .b (n_128), .cin (n_121));
FA__1_498 F41 (.carry (n_76), .sum (Result[9]), .a (n_75), .b (n_63), .cin (n_65));
FA__1_501 F33 (.carry (n_74), .sum (n_75), .a (n_73), .b (n_61), .cin (n_59));
FA__1_504 F29 (.carry (n_72), .sum (n_73), .a (n_69), .b (n_57), .cin (n_71));
FA__1_507 F24 (.carry (n_70), .sum (n_71), .a (n_119), .b (n_165), .cin (n_110));
FA__1_510 F18 (.carry (n_68), .sum (n_69), .a (n_67), .b (n_53), .cin (n_55));
FA__1_513 F6 (.carry (n_66), .sum (n_67), .a (n_143), .b (n_135), .cin (n_127));
FA__1_516 F40 (.carry (n_65), .sum (Result[8]), .a (n_64), .b (n_50), .cin (n_52));
FA__1_519 F32 (.carry (n_63), .sum (n_64), .a (n_62), .b (n_48), .cin (n_46));
FA__1_522 F28 (.carry (n_61), .sum (n_62), .a (n_58), .b (n_44), .cin (n_60));
FA__1_525 F23 (.carry (n_59), .sum (n_60), .a (n_42), .b (n_164), .cin (n_109));
FA__1_528 F17 (.carry (n_57), .sum (n_58), .a (n_54), .b (n_40), .cin (n_56));
FA__1_531 F10 (.carry (n_55), .sum (n_56), .a (n_134), .b (n_126), .cin (n_120));
HA__1_534 H1 (.c (n_53), .s (n_54), .a (n_150), .b (n_142));
FA__1_537 F39 (.carry (n_52), .sum (Result[7]), .a (n_51), .b (n_37), .cin (n_39));
FA__1_540 F31 (.carry (n_50), .sum (n_51), .a (n_49), .b (n_35), .cin (n_33));
FA__1_543 F27 (.carry (n_48), .sum (n_49), .a (n_45), .b (n_31), .cin (n_47));
FA__1_546 F22 (.carry (n_46), .sum (n_47), .a (n_29), .b (n_163), .cin (n_108));
FA__1_549 F16 (.carry (n_44), .sum (n_45), .a (n_41), .b (n_27), .cin (n_43));
FA__1_552 F9 (.carry (n_42), .sum (n_43), .a (n_133), .b (n_125), .cin (n_118));
FA__1_555 F5 (.carry (n_40), .sum (n_41), .a (n_157), .b (n_149), .cin (n_141));
FA__1_558 F38 (.carry (n_39), .sum (Result[6]), .a (n_38), .b (n_20), .cin (n_26));
HA__1_561 H13 (.c (n_37), .s (n_38), .a (n_36), .b (n_12));
FA__1_564 F26 (.carry (n_35), .sum (n_36), .a (n_32), .b (n_4), .cin (n_34));
HA__1_567 H6 (.c (n_33), .s (n_34), .a (n_162), .b (n_2));
FA__1_570 F15 (.carry (n_31), .sum (n_32), .a (n_28), .b (C), .cin (n_30));
FA__1_573 F8 (.carry (n_29), .sum (n_30), .a (n_132), .b (n_124), .cin (n_117));
FA__1_576 F4 (.carry (n_27), .sum (n_28), .a (n_156), .b (n_148), .cin (n_140));
HA__1_579 H15 (.c (n_26), .s (Result[5]), .a (n_21), .b (n_25));
HA__1_582 H11 (.c (n_25), .s (Result[4]), .a (n_19), .b (n_24));
HA__1_585 H7 (.c (n_24), .s (Result[3]), .a (n_17), .b (n_23));
HA__1_588 H4 (.c (n_23), .s (Result[2]), .a (n_15), .b (n_22));
HA__1_591 H0 (.c (n_22), .s (Result[1]), .a (n_158), .b (n_151));
HA__1_594 H12 (.c (n_20), .s (n_21), .a (n_13), .b (n_18));
HA__1_597 H8 (.c (n_18), .s (n_19), .a (n_11), .b (n_16));
FA__1_600 F12 (.carry (n_16), .sum (n_17), .a (n_7), .b (n_14), .cin (n_137));
FA__1_603 F0 (.carry (n_14), .sum (n_15), .a (n_159), .b (n_152), .cin (n_144));
FA__1_606 F25 (.carry (n_12), .sum (n_13), .a (n_5), .b (n_10), .cin (n_8));
FA__1_609 F13 (.carry (n_10), .sum (n_11), .a (n_1), .b (n_6), .cin (n_9));
HA__1_612 H2 (.c (n_8), .s (n_9), .a (n_138), .b (n_130));
FA__1_615 F1 (.carry (n_6), .sum (n_7), .a (n_160), .b (n_153), .cin (n_145));
FA__1_618 F14 (.carry (n_4), .sum (n_5), .a (S), .b (n_0), .cin (n_3));
FA__1_621 F7 (.carry (n_2), .sum (n_3), .a (n_131), .b (n_123), .cin (n_116));
FA__1_624 F2 (.carry (n_0), .sum (n_1), .a (n_161), .b (n_154), .cin (n_146));
FA__1_627 F3 (.carry (C), .sum (S), .a (n_155), .b (n_147), .cin (n_139));

endmodule //WTM8__1_628

module WTM32 (A, B, Result);

output [63:0] Result;
input [31:0] A;
input [31:0] B;
wire \P[0][15] ;
wire \P[0][14] ;
wire \P[0][13] ;
wire \P[0][12] ;
wire \P[0][11] ;
wire \P[0][10] ;
wire \P[0][9] ;
wire \P[0][8] ;
wire \P[0][7] ;
wire \P[0][6] ;
wire \P[0][5] ;
wire \P[0][4] ;
wire \P[0][3] ;
wire \P[0][2] ;
wire \P[0][1] ;
wire \couple[0][24] ;
wire \couple[0][23] ;
wire \couple[0][22] ;
wire \couple[0][21] ;
wire \couple[0][20] ;
wire \couple[0][19] ;
wire \couple[0][18] ;
wire \couple[0][17] ;
wire \couple[0][16] ;
wire \couple[0][15] ;
wire \couple[0][14] ;
wire \couple[0][13] ;
wire \couple[0][12] ;
wire \couple[0][11] ;
wire \couple[0][10] ;
wire \couple[0][9] ;
wire \couple[0][8] ;
wire \P[2][15] ;
wire \P[2][14] ;
wire \P[2][13] ;
wire \P[2][12] ;
wire \P[2][11] ;
wire \P[2][10] ;
wire \P[2][9] ;
wire \P[2][8] ;
wire \P[2][7] ;
wire \P[2][6] ;
wire \P[2][5] ;
wire \P[2][4] ;
wire \P[2][3] ;
wire \P[2][2] ;
wire \P[2][1] ;
wire \P[2][0] ;
wire \P[3][15] ;
wire \P[3][14] ;
wire \P[3][13] ;
wire \P[3][12] ;
wire \P[3][11] ;
wire \P[3][10] ;
wire \P[3][9] ;
wire \P[3][8] ;
wire \P[3][7] ;
wire \P[3][6] ;
wire \P[3][5] ;
wire \P[3][4] ;
wire \P[3][3] ;
wire \P[3][2] ;
wire \P[3][1] ;
wire \P[3][0] ;
wire \couple[1][40] ;
wire \couple[1][39] ;
wire \couple[1][38] ;
wire \couple[1][37] ;
wire \couple[1][36] ;
wire \couple[1][35] ;
wire \couple[1][34] ;
wire \couple[1][33] ;
wire \couple[1][32] ;
wire \couple[1][31] ;
wire \couple[1][30] ;
wire \couple[1][29] ;
wire \couple[1][28] ;
wire \couple[1][27] ;
wire \couple[1][26] ;
wire \couple[1][25] ;
wire \couple[1][24] ;
wire \Quadruple[0][41] ;
wire \Quadruple[0][40] ;
wire \Quadruple[0][39] ;
wire \Quadruple[0][38] ;
wire \Quadruple[0][37] ;
wire \Quadruple[0][36] ;
wire \Quadruple[0][35] ;
wire \Quadruple[0][34] ;
wire \Quadruple[0][33] ;
wire \Quadruple[0][32] ;
wire \Quadruple[0][31] ;
wire \Quadruple[0][30] ;
wire \Quadruple[0][29] ;
wire \Quadruple[0][28] ;
wire \Quadruple[0][27] ;
wire \Quadruple[0][26] ;
wire \Quadruple[0][25] ;
wire \Quadruple[0][24] ;
wire \Quadruple[0][23] ;
wire \Quadruple[0][22] ;
wire \Quadruple[0][21] ;
wire \Quadruple[0][20] ;
wire \Quadruple[0][19] ;
wire \Quadruple[0][18] ;
wire \Quadruple[0][17] ;
wire \Quadruple[0][16] ;
wire \P[4][15] ;
wire \P[4][14] ;
wire \P[4][13] ;
wire \P[4][12] ;
wire \P[4][11] ;
wire \P[4][10] ;
wire \P[4][9] ;
wire \P[4][8] ;
wire \P[4][7] ;
wire \P[4][6] ;
wire \P[4][5] ;
wire \P[4][4] ;
wire \P[4][3] ;
wire \P[4][2] ;
wire \P[4][1] ;
wire \P[4][0] ;
wire \P[5][15] ;
wire \P[5][14] ;
wire \P[5][13] ;
wire \P[5][12] ;
wire \P[5][11] ;
wire \P[5][10] ;
wire \P[5][9] ;
wire \P[5][8] ;
wire \P[5][7] ;
wire \P[5][6] ;
wire \P[5][5] ;
wire \P[5][4] ;
wire \P[5][3] ;
wire \P[5][2] ;
wire \P[5][1] ;
wire \P[5][0] ;
wire \couple[2][32] ;
wire \couple[2][31] ;
wire \couple[2][30] ;
wire \couple[2][29] ;
wire \couple[2][28] ;
wire \couple[2][27] ;
wire \couple[2][26] ;
wire \couple[2][25] ;
wire \couple[2][24] ;
wire \couple[2][23] ;
wire \couple[2][22] ;
wire \couple[2][21] ;
wire \couple[2][20] ;
wire \couple[2][19] ;
wire \couple[2][18] ;
wire \couple[2][17] ;
wire \couple[2][16] ;
wire \P[6][15] ;
wire \P[6][14] ;
wire \P[6][13] ;
wire \P[6][12] ;
wire \P[6][11] ;
wire \P[6][10] ;
wire \P[6][9] ;
wire \P[6][8] ;
wire \P[6][7] ;
wire \P[6][6] ;
wire \P[6][5] ;
wire \P[6][4] ;
wire \P[6][3] ;
wire \P[6][2] ;
wire \P[6][1] ;
wire \P[6][0] ;
wire \P[7][15] ;
wire \P[7][14] ;
wire \P[7][13] ;
wire \P[7][12] ;
wire \P[7][11] ;
wire \P[7][10] ;
wire \P[7][9] ;
wire \P[7][8] ;
wire \P[7][7] ;
wire \P[7][6] ;
wire \P[7][5] ;
wire \P[7][4] ;
wire \P[7][3] ;
wire \P[7][2] ;
wire \P[7][1] ;
wire \P[7][0] ;
wire \couple[3][48] ;
wire \couple[3][47] ;
wire \couple[3][46] ;
wire \couple[3][45] ;
wire \couple[3][44] ;
wire \couple[3][43] ;
wire \couple[3][42] ;
wire \couple[3][41] ;
wire \couple[3][40] ;
wire \couple[3][39] ;
wire \couple[3][38] ;
wire \couple[3][37] ;
wire \couple[3][36] ;
wire \couple[3][35] ;
wire \couple[3][34] ;
wire \couple[3][33] ;
wire \couple[3][32] ;
wire \Quadruple[1][49] ;
wire \Quadruple[1][48] ;
wire \Quadruple[1][47] ;
wire \Quadruple[1][46] ;
wire \Quadruple[1][45] ;
wire \Quadruple[1][44] ;
wire \Quadruple[1][43] ;
wire \Quadruple[1][42] ;
wire \Quadruple[1][41] ;
wire \Quadruple[1][40] ;
wire \Quadruple[1][39] ;
wire \Quadruple[1][38] ;
wire \Quadruple[1][37] ;
wire \Quadruple[1][36] ;
wire \Quadruple[1][35] ;
wire \Quadruple[1][34] ;
wire \Quadruple[1][33] ;
wire \Quadruple[1][32] ;
wire \Quadruple[1][31] ;
wire \Quadruple[1][30] ;
wire \Quadruple[1][29] ;
wire \Quadruple[1][28] ;
wire \Quadruple[1][27] ;
wire \Quadruple[1][26] ;
wire \Quadruple[1][25] ;
wire \Quadruple[1][24] ;
wire \Eight[0][50] ;
wire \Eight[0][49] ;
wire \Eight[0][48] ;
wire \Eight[0][47] ;
wire \Eight[0][46] ;
wire \Eight[0][45] ;
wire \Eight[0][44] ;
wire \Eight[0][43] ;
wire \Eight[0][42] ;
wire \Eight[0][41] ;
wire \Eight[0][40] ;
wire \Eight[0][39] ;
wire \Eight[0][38] ;
wire \Eight[0][37] ;
wire \Eight[0][36] ;
wire \Eight[0][35] ;
wire \Eight[0][34] ;
wire \Eight[0][33] ;
wire \Eight[0][32] ;
wire \Eight[0][31] ;
wire \Eight[0][30] ;
wire \Eight[0][29] ;
wire \Eight[0][28] ;
wire \Eight[0][27] ;
wire \Eight[0][26] ;
wire \Eight[0][25] ;
wire \Eight[0][24] ;
wire \Eight[0][23] ;
wire \Eight[0][22] ;
wire \Eight[0][21] ;
wire \Eight[0][20] ;
wire \Eight[0][19] ;
wire \Eight[0][18] ;
wire \Eight[0][17] ;
wire \Eight[0][16] ;
wire \Eight[0][15] ;
wire \Eight[0][14] ;
wire \Eight[0][13] ;
wire \Eight[0][12] ;
wire \Eight[0][11] ;
wire \Eight[0][10] ;
wire \Eight[0][9] ;
wire \Eight[0][8] ;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire \P[10][15] ;
wire \P[10][14] ;
wire \P[10][13] ;
wire \P[10][12] ;
wire \P[10][11] ;
wire \P[10][10] ;
wire \P[10][9] ;
wire \P[10][8] ;
wire \P[10][7] ;
wire \P[10][6] ;
wire \P[10][5] ;
wire \P[10][4] ;
wire \P[10][3] ;
wire \P[10][2] ;
wire \P[10][1] ;
wire \P[10][0] ;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_62;
wire \out[63] ;
wire \out[62] ;
wire \out[61] ;
wire \out[60] ;
wire \out[59] ;
wire \out[58] ;
wire \out[57] ;
wire \out[56] ;
wire \out[55] ;
wire \out[54] ;
wire \out[53] ;
wire \out[52] ;
wire \out[51] ;
wire \out[50] ;
wire \out[49] ;
wire \out[48] ;
wire \out[47] ;
wire \out[46] ;
wire \out[45] ;
wire \out[44] ;
wire \out[43] ;
wire \out[42] ;
wire \out[41] ;
wire \out[40] ;
wire \out[39] ;
wire \out[38] ;
wire \out[37] ;
wire \out[36] ;
wire \out[35] ;
wire \out[34] ;
wire \out[33] ;
wire \out[32] ;
wire \out[31] ;
wire \out[30] ;
wire \out[29] ;
wire \out[28] ;
wire \out[27] ;
wire \out[26] ;
wire \out[25] ;
wire \out[24] ;
wire \out[23] ;
wire \out[22] ;
wire \out[21] ;
wire \out[20] ;
wire \out[19] ;
wire \out[18] ;
wire \out[17] ;
wire \out[16] ;
wire \P[14][15] ;
wire \P[14][14] ;
wire \P[14][13] ;
wire \P[14][12] ;
wire \P[14][11] ;
wire \P[14][10] ;
wire \P[14][9] ;
wire \P[14][8] ;
wire \P[14][7] ;
wire \P[14][6] ;
wire \P[14][5] ;
wire \P[14][4] ;
wire \P[14][3] ;
wire \P[14][2] ;
wire \P[14][1] ;
wire \P[14][0] ;
wire \b[31] ;
wire \b[30] ;
wire \b[29] ;
wire \b[28] ;
wire \b[27] ;
wire \b[26] ;
wire \b[25] ;
wire \b[24] ;
wire \b[23] ;
wire \b[22] ;
wire \b[21] ;
wire \b[20] ;
wire \b[19] ;
wire \b[18] ;
wire \b[17] ;
wire \b[16] ;
wire \b[15] ;
wire \b[14] ;
wire \b[13] ;
wire \b[12] ;
wire \b[11] ;
wire \b[10] ;
wire \b[9] ;
wire \b[8] ;
wire \b[7] ;
wire \b[6] ;
wire \b[5] ;
wire \b[4] ;
wire \b[3] ;
wire \b[2] ;
wire \b[1] ;
wire \a[31] ;
wire \a[30] ;
wire \a[29] ;
wire \a[28] ;
wire \a[27] ;
wire \a[26] ;
wire \a[25] ;
wire \a[24] ;
wire \a[23] ;
wire \a[22] ;
wire \a[21] ;
wire \a[20] ;
wire \a[19] ;
wire \a[18] ;
wire \a[17] ;
wire \a[16] ;
wire \a[15] ;
wire \a[14] ;
wire \a[13] ;
wire \a[12] ;
wire \a[11] ;
wire \a[10] ;
wire \a[9] ;
wire \a[8] ;
wire \a[7] ;
wire \a[6] ;
wire \a[5] ;
wire \a[4] ;
wire \a[3] ;
wire \a[2] ;
wire \a[1] ;
wire n_0_0_0;
wire \couple[6][48] ;
wire \couple[6][47] ;
wire \couple[6][46] ;
wire \couple[6][45] ;
wire \couple[6][44] ;
wire \couple[6][43] ;
wire \couple[6][42] ;
wire \couple[6][41] ;
wire \couple[6][40] ;
wire \couple[6][39] ;
wire \couple[6][38] ;
wire \couple[6][37] ;
wire \couple[6][36] ;
wire \couple[6][35] ;
wire \couple[6][34] ;
wire \couple[6][33] ;
wire \couple[6][32] ;
wire \P[13][15] ;
wire \P[13][14] ;
wire \P[13][13] ;
wire \P[13][12] ;
wire \P[13][11] ;
wire \P[13][10] ;
wire \P[13][9] ;
wire \P[13][8] ;
wire \P[13][7] ;
wire \P[13][6] ;
wire \P[13][5] ;
wire \P[13][4] ;
wire \P[13][3] ;
wire \P[13][2] ;
wire \P[13][1] ;
wire \P[13][0] ;
wire \P[15][15] ;
wire \P[15][14] ;
wire \P[15][13] ;
wire \P[15][12] ;
wire \P[15][11] ;
wire \P[15][10] ;
wire \P[15][9] ;
wire \P[15][8] ;
wire \P[15][7] ;
wire \P[15][6] ;
wire \P[15][5] ;
wire \P[15][4] ;
wire \P[15][3] ;
wire \P[15][2] ;
wire \P[15][1] ;
wire \P[15][0] ;
wire \couple[7][63] ;
wire \couple[7][62] ;
wire \couple[7][61] ;
wire \couple[7][60] ;
wire \couple[7][59] ;
wire \couple[7][58] ;
wire \couple[7][57] ;
wire \couple[7][56] ;
wire \couple[7][55] ;
wire \couple[7][54] ;
wire \couple[7][53] ;
wire \couple[7][52] ;
wire \couple[7][51] ;
wire \couple[7][50] ;
wire \couple[7][49] ;
wire \couple[7][48] ;
wire \Quadruple[3][63] ;
wire \Quadruple[3][62] ;
wire \Quadruple[3][61] ;
wire \Quadruple[3][60] ;
wire \Quadruple[3][59] ;
wire \Quadruple[3][58] ;
wire \Quadruple[3][57] ;
wire \Quadruple[3][56] ;
wire \Quadruple[3][55] ;
wire \Quadruple[3][54] ;
wire \Quadruple[3][53] ;
wire \Quadruple[3][52] ;
wire \Quadruple[3][51] ;
wire \Quadruple[3][50] ;
wire \Quadruple[3][49] ;
wire \Quadruple[3][48] ;
wire \Quadruple[3][47] ;
wire \Quadruple[3][46] ;
wire \Quadruple[3][45] ;
wire \Quadruple[3][44] ;
wire \Quadruple[3][43] ;
wire \Quadruple[3][42] ;
wire \Quadruple[3][41] ;
wire \Quadruple[3][40] ;
wire \Eight[1][63] ;
wire \Eight[1][62] ;
wire \Eight[1][61] ;
wire \Eight[1][60] ;
wire \Eight[1][59] ;
wire \Eight[1][58] ;
wire \Eight[1][57] ;
wire \Eight[1][56] ;
wire \Eight[1][55] ;
wire \Eight[1][54] ;
wire \Eight[1][53] ;
wire \Eight[1][52] ;
wire \Eight[1][51] ;
wire \Eight[1][50] ;
wire \Eight[1][49] ;
wire \Eight[1][48] ;
wire \Eight[1][47] ;
wire \Eight[1][46] ;
wire \Eight[1][45] ;
wire \Eight[1][44] ;
wire \Eight[1][43] ;
wire \Eight[1][42] ;
wire \Eight[1][41] ;
wire \Eight[1][40] ;
wire \Eight[1][39] ;
wire \Eight[1][38] ;
wire \Eight[1][37] ;
wire \Eight[1][36] ;
wire \Eight[1][35] ;
wire \Eight[1][34] ;
wire \Eight[1][33] ;
wire \Eight[1][32] ;
wire \Eight[1][31] ;
wire \Eight[1][30] ;
wire \Eight[1][29] ;
wire \Eight[1][28] ;
wire \Eight[1][27] ;
wire \Eight[1][26] ;
wire \Eight[1][25] ;
wire \Eight[1][24] ;
wire \Eight[1][23] ;
wire \Eight[1][22] ;
wire \Eight[1][21] ;
wire \Eight[1][20] ;
wire \Eight[1][19] ;
wire \Eight[1][18] ;
wire \Eight[1][17] ;
wire \Eight[1][16] ;
wire \P[12][15] ;
wire \P[12][14] ;
wire \P[12][13] ;
wire \P[12][12] ;
wire \P[12][11] ;
wire \P[12][10] ;
wire \P[12][9] ;
wire \P[12][8] ;
wire \P[12][7] ;
wire \P[12][6] ;
wire \P[12][5] ;
wire \P[12][4] ;
wire \P[12][3] ;
wire \P[12][2] ;
wire \P[12][1] ;
wire \P[12][0] ;
wire \Quadruple[2][57] ;
wire \Quadruple[2][56] ;
wire \Quadruple[2][55] ;
wire \Quadruple[2][54] ;
wire \Quadruple[2][53] ;
wire \Quadruple[2][52] ;
wire \Quadruple[2][51] ;
wire \Quadruple[2][50] ;
wire \Quadruple[2][49] ;
wire \Quadruple[2][48] ;
wire \Quadruple[2][47] ;
wire \Quadruple[2][46] ;
wire \Quadruple[2][45] ;
wire \Quadruple[2][44] ;
wire \Quadruple[2][43] ;
wire \Quadruple[2][42] ;
wire \Quadruple[2][41] ;
wire \Quadruple[2][40] ;
wire \Quadruple[2][39] ;
wire \Quadruple[2][38] ;
wire \Quadruple[2][37] ;
wire \Quadruple[2][36] ;
wire \Quadruple[2][35] ;
wire \Quadruple[2][34] ;
wire \Quadruple[2][33] ;
wire \Quadruple[2][32] ;
wire \couple[5][56] ;
wire \couple[5][55] ;
wire \couple[5][54] ;
wire \couple[5][53] ;
wire \couple[5][52] ;
wire \couple[5][51] ;
wire \couple[5][50] ;
wire \couple[5][49] ;
wire \couple[5][48] ;
wire \couple[5][47] ;
wire \couple[5][46] ;
wire \couple[5][45] ;
wire \couple[5][44] ;
wire \couple[5][43] ;
wire \couple[5][42] ;
wire \couple[5][41] ;
wire \couple[5][40] ;
wire \P[11][15] ;
wire \P[11][14] ;
wire \P[11][13] ;
wire \P[11][12] ;
wire \P[11][11] ;
wire \P[11][10] ;
wire \P[11][9] ;
wire \P[11][8] ;
wire \P[11][7] ;
wire \P[11][6] ;
wire \P[11][5] ;
wire \P[11][4] ;
wire \P[11][3] ;
wire \P[11][2] ;
wire \P[11][1] ;
wire \P[11][0] ;
wire spw__n325;
wire spw__n324;
wire spw__n278;
wire spw__n277;
wire spw__n276;
wire spw__n314;
wire spw__n230;
wire spw__n229;
wire spw__n228;
wire spw__n227;
wire spw__n226;
wire spw__n225;
wire spw__n216;
wire spw__n215;
wire spw__n184;
wire spw__n183;
wire spw__n182;
wire spw__n167;
wire spw__n166;
wire spw__n155;
wire \couple[4][40] ;
wire \couple[4][39] ;
wire \couple[4][38] ;
wire \couple[4][37] ;
wire \couple[4][36] ;
wire \couple[4][35] ;
wire \couple[4][34] ;
wire \couple[4][33] ;
wire \couple[4][32] ;
wire \couple[4][31] ;
wire \couple[4][30] ;
wire \couple[4][29] ;
wire \couple[4][28] ;
wire \couple[4][27] ;
wire \couple[4][26] ;
wire \couple[4][25] ;
wire \couple[4][24] ;
wire spw__n154;
wire spw__n153;
wire spw__n152;
wire spw__n139;
wire spw__n138;
wire spw__n137;
wire spw__n136;
wire spw__n135;
wire spw__n124;
wire spw__n123;
wire spw__n122;
wire spw__n113;
wire spw__n112;
wire spw__n111;
wire spw__n90;
wire spw__n89;
wire spw__n88;
wire spw__n81;
wire spw__n80;
wire spw__n384;
wire spw__n67;
wire spw__n54;
wire spw__n53;
wire \P[9][15] ;
wire \P[9][14] ;
wire \P[9][13] ;
wire \P[9][12] ;
wire \P[9][11] ;
wire \P[9][10] ;
wire \P[9][9] ;
wire \P[9][8] ;
wire \P[9][7] ;
wire \P[9][6] ;
wire \P[9][5] ;
wire \P[9][4] ;
wire \P[9][3] ;
wire \P[9][2] ;
wire \P[9][1] ;
wire \P[9][0] ;
wire \P[8][15] ;
wire \P[8][14] ;
wire \P[8][13] ;
wire \P[8][12] ;
wire \P[8][11] ;
wire \P[8][10] ;
wire \P[8][9] ;
wire \P[8][8] ;
wire spw__n52;
wire spw__n51;
wire spw__n50;
wire spt__n12;
wire spt__n9;
wire spt__n6;
wire spt__n3;
wire sps__n1;
wire \P[1][15] ;
wire \P[1][14] ;
wire \P[1][13] ;
wire \P[1][12] ;
wire \P[1][11] ;
wire \P[1][10] ;
wire \P[1][9] ;
wire \P[1][8] ;
wire \P[1][7] ;
wire \P[1][6] ;
wire \P[1][5] ;
wire \P[1][4] ;
wire \P[1][3] ;
wire \P[1][2] ;
wire \P[1][1] ;
wire \P[1][0] ;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire uc_65;
wire uc_66;
wire uc_67;
wire uc_68;
wire uc_69;
wire uc_70;
wire uc_71;
wire uc_72;
wire uc_73;
wire uc_74;
wire uc_75;
wire uc_76;
wire uc_77;
wire uc_78;
wire uc_79;
wire uc_80;
wire uc_81;
wire uc_82;
wire uc_83;
wire uc_84;
wire uc_85;
wire uc_86;
wire uc_87;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;
wire uc_94;
wire uc_95;
wire uc_96;
wire uc_97;
wire uc_98;
wire uc_99;
wire uc_100;
wire uc_101;
wire uc_102;
wire uc_103;
wire uc_104;
wire uc_105;
wire uc_106;
wire uc_107;
wire uc_108;
wire uc_109;
wire uc_110;
wire uc_111;
wire uc_112;
wire uc_113;
wire uc_114;
wire uc_115;
wire uc_116;
wire uc_117;
wire uc_118;
wire uc_119;
wire uc_120;
wire uc_121;
wire uc_122;
wire uc_123;
wire uc_124;
wire uc_125;
wire uc_126;
wire uc_127;
wire uc_128;
wire uc_129;
wire uc_130;
wire uc_131;
wire uc_132;
wire uc_133;
wire uc_134;
wire uc_135;
wire uc_136;
wire uc_137;
wire uc_138;
wire uc_139;
wire uc_140;
wire uc_141;
wire uc_142;
wire uc_143;
wire uc_144;
wire uc_145;
wire uc_146;
wire uc_147;
wire uc_148;
wire uc_149;
wire uc_150;
wire uc_151;
wire uc_152;
wire uc_153;
wire uc_154;
wire uc_155;
wire uc_156;
wire uc_157;
wire uc_158;
wire uc_159;
wire uc_160;
wire uc_161;
wire uc_162;
wire uc_163;
wire uc_164;
wire uc_165;
wire uc_166;
wire uc_167;
wire uc_168;
wire uc_169;
wire uc_170;
wire uc_171;
wire uc_172;
wire uc_173;
wire uc_174;
wire uc_175;
wire uc_176;
wire uc_177;
wire uc_178;
wire uc_179;
wire uc_180;
wire uc_181;
wire uc_182;
wire uc_183;
wire uc_184;
wire uc_185;
wire uc_186;
wire uc_187;
wire uc_188;
wire uc_189;
wire uc_190;
wire uc_191;
wire uc_192;
wire uc_193;
wire uc_194;
wire uc_195;
wire uc_196;
wire uc_197;
wire uc_198;
wire uc_199;
wire uc_200;
wire uc_201;
wire uc_202;
wire uc_203;
wire uc_204;
wire uc_205;
wire uc_206;
wire uc_207;
wire uc_208;
wire uc_209;
wire uc_210;
wire uc_211;
wire uc_212;
wire uc_213;
wire uc_214;
wire uc_215;
wire uc_216;
wire uc_217;
wire uc_218;
wire uc_219;
wire uc_220;
wire uc_221;
wire uc_222;
wire uc_223;
wire uc_224;
wire uc_225;
wire uc_226;
wire uc_227;
wire uc_228;
wire uc_229;
wire uc_230;
wire uc_231;
wire uc_232;
wire uc_233;
wire uc_234;
wire uc_235;
wire uc_236;
wire uc_237;
wire uc_238;
wire uc_239;
wire uc_240;
wire uc_241;
wire uc_242;
wire uc_243;
wire uc_244;
wire uc_245;
wire uc_246;
wire uc_247;
wire uc_248;
wire uc_249;
wire uc_250;
wire uc_251;
wire uc_252;
wire uc_253;
wire uc_254;
wire uc_255;
wire uc_256;
wire uc_257;
wire uc_258;
wire uc_259;
wire uc_260;
wire uc_261;
wire uc_262;
wire uc_263;
wire uc_264;
wire uc_265;
wire uc_266;
wire uc_267;
wire uc_268;
wire uc_269;
wire uc_270;
wire uc_271;
wire uc_272;
wire uc_273;
wire uc_274;
wire uc_275;
wire uc_276;
wire uc_277;
wire uc_278;
wire uc_279;
wire uc_280;
wire uc_281;
wire uc_282;
wire uc_283;
wire uc_284;
wire uc_285;
wire uc_286;
wire uc_287;
wire uc_288;
wire uc_289;
wire uc_290;
wire uc_291;
wire uc_292;
wire uc_293;
wire uc_294;
wire uc_295;
wire uc_296;
wire uc_297;
wire uc_298;
wire uc_299;
wire uc_300;
wire uc_301;
wire uc_302;
wire uc_303;
wire uc_304;
wire uc_305;
wire uc_306;
wire uc_307;
wire uc_308;
wire uc_309;
wire uc_310;
wire uc_311;
wire uc_312;
wire uc_313;
wire uc_314;
wire uc_315;
wire uc_316;
wire uc_317;
wire uc_318;
wire uc_319;
wire uc_320;
wire uc_321;
wire uc_322;
wire uc_323;
wire uc_324;
wire uc_325;
wire uc_326;
wire uc_327;
wire uc_328;
wire uc_329;
wire uc_330;
wire uc_331;
wire uc_332;
wire uc_333;
wire uc_334;
wire uc_335;
wire uc_336;
wire uc_337;
wire uc_338;
wire uc_339;
wire uc_340;
wire uc_341;
wire uc_342;
wire uc_343;
wire uc_344;
wire uc_345;
wire uc_346;
wire uc_347;
wire uc_348;
wire uc_349;
wire uc_350;
wire uc_351;
wire uc_352;
wire uc_353;
wire uc_354;
wire uc_355;
wire uc_356;
wire uc_357;
wire uc_358;
wire uc_359;
wire uc_360;
wire uc_361;
wire uc_362;
wire uc_363;
wire uc_364;
wire uc_365;
wire uc_366;
wire uc_367;
wire uc_368;
wire uc_369;
wire uc_370;
wire uc_371;
wire uc_372;
wire uc_373;
wire uc_374;
wire uc_375;
wire uc_376;
wire uc_377;
wire uc_378;
wire uc_379;
wire uc_380;
wire uc_381;
wire uc_382;
wire uc_383;
wire uc_384;
wire uc_385;
wire uc_386;
wire uc_387;
wire uc_388;
wire uc_389;
wire uc_390;
wire uc_391;
wire uc_392;
wire uc_393;
wire uc_394;
wire uc_395;
wire uc_396;
wire uc_397;
wire uc_398;
wire uc_399;
wire uc_400;
wire uc_401;
wire uc_402;
wire uc_403;
wire uc_404;
wire uc_405;
wire uc_406;
wire uc_407;
wire uc_408;
wire uc_409;
wire uc_410;
wire uc_411;
wire uc_412;
wire uc_413;
wire uc_414;
wire uc_415;
wire uc_416;
wire uc_417;
wire uc_418;
wire uc_419;
wire uc_420;
wire uc_421;
wire uc_422;
wire uc_423;
wire uc_424;
wire uc_425;
wire uc_426;
wire uc_427;
wire uc_428;
wire uc_429;
wire uc_430;
wire uc_431;
wire uc_432;
wire uc_433;
wire uc_434;
wire uc_435;
wire uc_436;
wire uc_437;
wire uc_438;
wire uc_439;
wire uc_440;
wire uc_441;
wire uc_442;
wire uc_443;
wire uc_444;
wire uc_445;
wire uc_446;
wire uc_447;
wire uc_448;
wire uc_449;
wire uc_450;
wire uc_451;
wire uc_452;
wire uc_453;
wire uc_454;
wire uc_455;
wire uc_456;
wire uc_457;
wire uc_458;
wire uc_459;
wire uc_460;
wire uc_461;
wire uc_462;
wire uc_463;
wire uc_464;
wire uc_465;
wire uc_466;
wire uc_467;
wire uc_468;
wire uc_469;
wire uc_470;
wire uc_471;
wire uc_472;
wire uc_473;
wire uc_474;
wire uc_475;
wire uc_476;
wire uc_477;
wire uc_478;
wire uc_479;
wire uc_480;
wire uc_481;
wire uc_482;
wire uc_483;
wire uc_484;
wire uc_485;
wire uc_486;
wire uc_487;
wire uc_488;
wire uc_489;
wire uc_490;
wire uc_491;
wire uc_492;
wire uc_493;
wire uc_494;
wire uc_495;
wire uc_496;
wire uc_497;
wire uc_498;
wire uc_499;
wire uc_500;
wire uc_501;
wire uc_502;
wire uc_503;
wire uc_504;
wire uc_505;
wire uc_506;
wire uc_507;
wire uc_508;
wire uc_509;
wire uc_510;
wire uc_511;
wire uc_512;
wire uc_513;
wire uc_514;
wire uc_515;
wire uc_516;
wire uc_517;
wire uc_518;
wire uc_519;
wire uc_520;
wire uc_521;
wire uc_522;
wire uc_523;
wire uc_524;
wire uc_525;
wire uc_526;
wire uc_527;
wire uc_528;
wire uc_529;
wire uc_530;
wire uc_531;
wire uc_532;
wire uc_533;
wire uc_534;
wire uc_535;
wire uc_536;
wire uc_537;
wire uc_538;
wire uc_539;
wire uc_540;
wire uc_541;
wire uc_542;
wire uc_543;
wire uc_544;
wire uc_545;
wire uc_546;
wire uc_547;
wire uc_548;
wire uc_549;
wire uc_550;
wire uc_551;
wire uc_552;
wire uc_553;
wire uc_554;
wire uc_555;
wire uc_556;
wire uc_557;
wire uc_558;
wire uc_559;
wire uc_560;
wire uc_561;
wire uc_562;
wire uc_563;
wire uc_564;
wire uc_565;
wire uc_566;
wire uc_567;
wire uc_568;
wire uc_569;
wire uc_570;
wire uc_571;
wire uc_572;
wire uc_573;
wire uc_574;
wire uc_575;
wire uc_576;
wire uc_577;
wire uc_578;
wire uc_579;
wire uc_580;
wire uc_581;
wire uc_582;
wire uc_583;
wire uc_584;
wire uc_585;
wire uc_586;
wire uc_587;
wire uc_588;
wire uc_589;
wire uc_590;
wire uc_591;
wire uc_592;
wire uc_593;
wire uc_594;
wire uc_595;
wire uc_596;
wire uc_597;
wire uc_598;
wire uc_599;
wire uc_600;
wire uc_601;
wire uc_602;
wire uc_603;
wire uc_604;
wire uc_605;
wire uc_606;
wire uc_607;
wire uc_608;
wire uc_609;
wire uc_610;
wire uc_611;
wire uc_612;
wire uc_613;
wire uc_614;
wire uc_615;
wire uc_616;
wire uc_617;
wire uc_618;
wire uc_619;
wire uc_620;
wire uc_621;
wire uc_622;
wire uc_623;
wire uc_624;
wire uc_625;
wire uc_626;
wire uc_627;
wire uc_628;
wire uc_629;
wire uc_630;
wire uc_631;
wire uc_632;
wire uc_633;
wire uc_634;
wire uc_635;
wire uc_636;
wire uc_637;
wire uc_638;
wire uc_639;
wire uc_640;
wire uc_641;
wire uc_642;
wire uc_643;
wire uc_644;
wire uc_645;
wire uc_646;
wire uc_647;
wire uc_648;
wire uc_649;
wire uc_650;
wire uc_651;
wire uc_652;
wire uc_653;
wire uc_654;
wire uc_655;
wire uc_656;
wire uc_657;
wire uc_658;
wire uc_659;
wire uc_660;
wire uc_661;
wire uc_662;
wire uc_663;
wire uc_664;
wire uc_665;
wire uc_666;
wire uc_667;
wire uc_668;
wire uc_669;
wire uc_670;
wire uc_671;
wire uc_672;
wire uc_673;
wire uc_674;
wire uc_675;
wire uc_676;
wire uc_677;
wire uc_678;
wire uc_679;
wire uc_680;
wire uc_681;
wire uc_682;
wire uc_683;
wire uc_684;
wire uc_685;
wire uc_686;
wire uc_687;
wire uc_688;
wire uc_689;
wire uc_690;
wire uc_691;
wire uc_692;
wire uc_693;
wire uc_694;
wire uc_695;
wire uc_696;
wire uc_697;
wire uc_698;
wire uc_699;
wire uc_700;
wire uc_701;
wire uc_702;
wire uc_703;
wire uc_704;
wire uc_705;
wire uc_706;
wire uc_707;
wire uc_708;
wire uc_709;
wire uc_710;
wire uc_711;
wire uc_712;
wire uc_713;
wire uc_714;
wire uc_715;
wire uc_716;
wire uc_717;
wire uc_718;
wire uc_719;
wire uc_720;
wire uc_721;
wire uc_722;
wire uc_723;
wire uc_724;
wire uc_725;
wire uc_726;
wire uc_727;
wire uc_728;
wire uc_729;
wire uc_730;
wire uc_731;
wire uc_732;
wire uc_733;
wire uc_734;
wire uc_735;
wire uc_736;
wire uc_737;
wire uc_738;
wire uc_739;
wire uc_740;
wire uc_741;
wire uc_742;
wire uc_743;
wire uc_744;
wire uc_745;
wire uc_746;
wire uc_747;
wire uc_748;
wire uc_749;
wire uc_750;
wire uc_751;
wire uc_752;
wire uc_753;
wire uc_754;
wire uc_755;
wire uc_756;
wire uc_757;
wire uc_758;
wire uc_759;
wire uc_760;
wire uc_761;
wire uc_762;
wire uc_763;
wire uc_764;
wire uc_765;
wire uc_766;
wire uc_767;
wire uc_768;
wire uc_769;
wire uc_770;
wire uc_771;
wire uc_772;
wire uc_773;
wire uc_774;
wire uc_775;
wire uc_776;
wire uc_777;
wire uc_778;
wire uc_779;
wire uc_780;
wire uc_781;
wire uc_782;
wire uc_783;
wire uc_784;
wire uc_785;
wire uc_786;
wire uc_787;
wire uc_788;
wire uc_789;
wire uc_790;
wire uc_791;
wire uc_792;
wire uc_793;
wire uc_794;
wire uc_795;
wire uc_796;
wire uc_797;
wire uc_798;
wire uc_799;
wire uc_800;
wire uc_801;
wire uc_802;
wire uc_803;
wire uc_804;
wire uc_805;
wire uc_806;
wire uc_807;
wire uc_808;
wire uc_809;
wire uc_810;
wire uc_811;
wire uc_812;
wire uc_813;
wire uc_814;
wire uc_815;
wire uc_816;
wire uc_817;
wire uc_818;
wire uc_819;
wire uc_820;
wire uc_821;
wire uc_822;
wire uc_823;
wire uc_824;
wire uc_825;
wire uc_826;
wire uc_827;
wire uc_828;
wire uc_829;
wire uc_830;
wire uc_831;
wire uc_832;
wire uc_833;
wire uc_834;
wire uc_835;
wire uc_836;
wire uc_837;
wire uc_838;
wire uc_839;
wire uc_840;
wire uc_841;
wire uc_842;
wire uc_843;
wire uc_844;
wire uc_845;
wire uc_846;
wire uc_847;
wire uc_848;
wire uc_849;
wire uc_850;
wire uc_851;
wire uc_852;
wire uc_853;
wire uc_854;
wire uc_855;
wire uc_856;
wire uc_857;
wire uc_858;
wire uc_859;
wire uc_860;
wire uc_861;
wire uc_862;
wire uc_863;
wire uc_864;
wire uc_865;
wire uc_866;
wire uc_867;
wire uc_868;
wire uc_869;
wire uc_870;
wire uc_871;
wire uc_872;
wire uc_873;
wire uc_874;
wire uc_875;
wire uc_876;
wire uc_877;
wire uc_878;
wire uc_879;
wire uc_880;
wire uc_881;
wire uc_882;
wire uc_883;
wire uc_884;
wire uc_885;
wire uc_886;
wire uc_887;
wire uc_888;
wire uc_889;
wire uc_890;
wire uc_891;
wire uc_892;
wire uc_893;
wire uc_894;
wire uc_895;
wire uc_896;
wire uc_897;
wire uc_898;
wire uc_899;
wire uc_900;
wire uc_901;
wire uc_902;
wire uc_903;
wire uc_904;
wire uc_905;
wire uc_906;
wire uc_907;
wire uc_908;
wire uc_909;
wire uc_910;
wire uc_911;
wire uc_912;
wire uc_913;
wire uc_914;
wire uc_915;
wire uc_916;
wire uc_917;
wire uc_918;
wire uc_919;
wire uc_920;
wire uc_921;
wire uc_922;
wire uc_923;
wire uc_924;
wire uc_925;
wire uc_926;
wire uc_927;
wire uc_928;
wire uc_929;
wire uc_930;
wire uc_931;
wire uc_932;
wire uc_933;
wire uc_934;
wire uc_935;
wire uc_936;
wire uc_937;
wire uc_938;
wire uc_939;
wire uc_940;
wire uc_941;
wire uc_942;
wire uc_943;
wire uc_944;
wire uc_945;
wire uc_946;
wire uc_947;
wire uc_948;
wire uc_949;
wire uc_950;
wire uc_951;
wire uc_952;
wire uc_953;
wire uc_954;
wire uc_955;
wire uc_956;
wire uc_957;
wire uc_958;
wire uc_959;
wire uc_960;
wire uc_961;
wire uc_962;
wire uc_963;
wire uc_964;
wire uc_965;
wire uc_966;
wire uc_967;
wire uc_968;
wire uc_969;
wire uc_970;
wire uc_971;
wire uc_972;
wire uc_973;
wire uc_974;
wire uc_975;
wire uc_976;
wire uc_977;
wire uc_978;
wire uc_979;
wire uc_980;
wire uc_981;
wire uc_982;
wire uc_983;
wire uc_984;
wire uc_985;
wire uc_986;
wire uc_987;
wire uc_988;
wire uc_989;
wire uc_990;
wire uc_991;
wire uc_992;
wire uc_993;
wire uc_994;
wire uc_995;
wire uc_996;
wire uc_997;
wire uc_998;
wire uc_999;
wire uc_1000;
wire uc_1001;
wire uc_1002;
wire uc_1003;
wire uc_1004;
wire uc_1005;
wire uc_1006;
wire uc_1007;
wire uc_1008;
wire uc_1009;
wire uc_1010;
wire uc_1011;
wire uc_1012;
wire uc_1013;
wire uc_1014;
wire uc_1015;
wire uc_1016;
wire uc_1017;
wire uc_1018;
wire uc_1019;
wire uc_1020;
wire uc_1021;
wire uc_1022;
wire uc_1023;
wire uc_1024;
wire uc_1025;
wire uc_1026;
wire uc_1027;
wire uc_1028;
wire uc_1029;
wire uc_1030;
wire uc_1031;
wire uc_1032;
wire uc_1033;
wire uc_1034;
wire uc_1035;
wire uc_1036;
wire uc_1037;
wire uc_1038;
wire uc_1039;
wire uc_1040;
wire uc_1041;
wire uc_1042;
wire uc_1043;
wire uc_1044;
wire uc_1045;
wire uc_1046;
wire uc_1047;
wire uc_1048;
wire uc_1049;
wire uc_1050;
wire uc_1051;
wire uc_1052;
wire uc_1053;
wire uc_1054;
wire uc_1055;
wire uc_1056;
wire uc_1057;
wire uc_1058;
wire uc_1059;
wire uc_1060;
wire uc_1061;
wire uc_1062;
wire uc_1063;
wire uc_1064;
wire uc_1065;
wire uc_1066;
wire uc_1067;
wire uc_1068;
wire uc_1069;
wire uc_1070;
wire uc_1071;
wire uc_1072;
wire uc_1073;
wire uc_1074;
wire uc_1075;
wire uc_1076;
wire uc_1077;
wire uc_1078;
wire uc_1079;
wire uc_1080;
wire uc_1081;
wire uc_1082;
wire uc_1083;
wire uc_1084;
wire uc_1085;
wire uc_1086;
wire uc_1087;
wire uc_1088;
wire uc_1089;
wire uc_1090;
wire uc_1091;
wire uc_1092;
wire uc_1093;
wire uc_1094;
wire uc_1095;
wire uc_1096;
wire uc_1097;
wire uc_1098;
wire uc_1099;
wire uc_1100;
wire uc_1101;
wire uc_1102;
wire uc_1103;
wire uc_1104;
wire uc_1105;
wire uc_1106;
wire uc_1107;
wire uc_1108;
wire uc_1109;
wire uc_1110;
wire uc_1111;
wire uc_1112;
wire uc_1113;
wire uc_1114;
wire uc_1115;
wire uc_1116;
wire uc_1117;
wire uc_1118;
wire uc_1119;
wire uc_1120;
wire uc_1121;
wire uc_1122;
wire uc_1123;
wire uc_1124;
wire uc_1125;
wire uc_1126;
wire uc_1127;
wire uc_1128;
wire uc_1129;
wire uc_1130;
wire uc_1131;
wire uc_1132;
wire uc_1133;
wire uc_1134;
wire uc_1135;
wire uc_1136;
wire uc_1137;
wire uc_1138;
wire uc_1139;
wire uc_1140;
wire uc_1141;
wire uc_1142;
wire uc_1143;
wire uc_1144;
wire uc_1145;
wire uc_1146;
wire uc_1147;
wire uc_1148;
wire uc_1149;
wire uc_1150;
wire uc_1151;
wire uc_1152;
wire uc_1153;
wire uc_1154;
wire uc_1155;
wire uc_1156;
wire uc_1157;
wire uc_1158;
wire uc_1159;
wire uc_1160;
wire uc_1161;
wire uc_1162;
wire uc_1163;
wire uc_1164;
wire uc_1165;
wire uc_1166;
wire uc_1167;
wire uc_1168;
wire uc_1169;
wire uc_1170;
wire uc_1171;
wire uc_1172;
wire uc_1173;
wire uc_1174;
wire uc_1175;
wire uc_1176;
wire uc_1177;
wire uc_1178;
wire uc_1179;
wire uc_1180;
wire uc_1181;
wire uc_1182;
wire uc_1183;
wire uc_1184;
wire uc_1185;
wire uc_1186;
wire uc_1187;
wire uc_1188;
wire uc_1189;
wire uc_1190;
wire uc_1191;
wire uc_1192;
wire uc_1193;
wire uc_1194;
wire uc_1195;
wire uc_1196;
wire uc_1197;
wire uc_1198;
wire uc_1199;
wire uc_1200;
wire uc_1201;
wire uc_1202;
wire uc_1203;
wire uc_1204;
wire uc_1205;
wire uc_1206;
wire uc_1207;
wire uc_1208;
wire uc_1209;
wire uc_1210;
wire uc_1211;
wire uc_1212;
wire uc_1213;
wire uc_1214;
wire uc_1215;
wire uc_1216;
wire uc_1217;
wire uc_1218;
wire uc_1219;
wire uc_1220;
wire uc_1221;
wire uc_1222;
wire uc_1223;
wire uc_1224;
wire uc_1225;
wire uc_1226;
wire uc_1227;
wire uc_1228;
wire uc_1229;
wire uc_1230;
wire uc_1231;
wire uc_1232;
wire uc_1233;
wire uc_1234;
wire uc_1235;
wire uc_1236;
wire uc_1237;
wire uc_1238;
wire uc_1239;
wire uc_1240;
wire uc_1241;
wire uc_1242;
wire uc_1243;
wire uc_1244;
wire uc_1245;
wire uc_1246;
wire uc_1247;
wire uc_1248;
wire uc_1249;
wire uc_1250;
wire uc_1251;
wire uc_1252;
wire uc_1253;
wire uc_1254;
wire uc_1255;
wire uc_1256;
wire uc_1257;
wire uc_1258;
wire uc_1259;
wire uc_1260;
wire uc_1261;
wire uc_1262;
wire uc_1263;
wire uc_1264;
wire uc_1265;
wire uc_1266;
wire uc_1267;
wire uc_1268;
wire uc_1269;
wire uc_1270;
wire uc_1271;
wire uc_1272;
wire uc_1273;
wire uc_1274;
wire uc_1275;
wire uc_1276;
wire uc_1277;
wire uc_1278;
wire uc_1279;
wire uc_1280;
wire uc_1281;
wire uc_1282;
wire uc_1283;
wire uc_1284;
wire uc_1285;
wire uc_1286;
wire uc_1287;
wire uc_1288;
wire uc_1289;
wire uc_1290;
wire uc_1291;
wire uc_1292;
wire uc_1293;
wire uc_1294;
wire uc_1295;
wire uc_1296;
wire uc_1297;
wire uc_1298;
wire uc_1299;
wire uc_1300;
wire uc_1301;
wire uc_1302;
wire uc_1303;
wire uc_1304;
wire uc_1305;
wire uc_1306;
wire uc_1307;
wire uc_1308;
wire uc_1309;
wire uc_1310;
wire uc_1311;
wire uc_1312;
wire uc_1313;
wire uc_1314;
wire uc_1315;
wire uc_1316;
wire uc_1317;
wire uc_1318;
wire uc_1319;
wire uc_1320;
wire uc_1321;
wire uc_1322;
wire uc_1323;
wire uc_1324;
wire uc_1325;
wire uc_1326;
wire uc_1327;
wire uc_1328;
wire uc_1329;
wire uc_1330;
wire uc_1331;
wire uc_1332;
wire uc_1333;
wire uc_1334;
wire uc_1335;
wire uc_1336;
wire uc_1337;
wire uc_1338;
wire uc_1339;
wire uc_1340;
wire uc_1341;
wire uc_1342;
wire uc_1343;
wire uc_1344;
wire uc_1345;
wire uc_1346;
wire uc_1347;
wire uc_1348;
wire uc_1349;
wire uc_1350;
wire uc_1351;
wire uc_1352;
wire uc_1353;
wire uc_1354;
wire uc_1355;
wire uc_1356;
wire uc_1357;
wire uc_1358;
wire uc_1359;
wire uc_1360;
wire uc_1361;
wire uc_1362;
wire uc_1363;
wire uc_1364;
wire uc_1365;
wire uc_1366;
wire uc_1367;
wire uc_1368;
wire uc_1369;
wire uc_1370;
wire uc_1371;
wire uc_1372;
wire uc_1373;
wire uc_1374;
wire uc_1375;
wire uc_1376;
wire uc_1377;
wire uc_1378;
wire uc_1379;
wire uc_1380;
wire uc_1381;
wire uc_1382;
wire uc_1383;
wire uc_1384;
wire uc_1385;
wire uc_1386;
wire uc_1387;
wire uc_1388;
wire uc_1389;
wire uc_1390;
wire uc_1391;
wire uc_1392;
wire uc_1393;
wire uc_1394;
wire uc_1395;
wire uc_1396;
wire uc_1397;
wire uc_1398;
wire uc_1399;
wire uc_1400;
wire uc_1401;
wire uc_1402;
wire uc_1403;
wire uc_1404;
wire uc_1405;
wire uc_1406;
wire uc_1407;
wire uc_1408;
wire uc_1409;
wire uc_1410;
wire uc_1411;
wire uc_1412;
wire uc_1413;
wire uc_1414;
wire uc_1415;
wire uc_1416;
wire uc_1417;
wire uc_1418;
wire uc_1419;
wire uc_1420;
wire uc_1421;
wire uc_1422;
wire uc_1423;
wire uc_1424;
wire uc_1425;
wire uc_1426;
wire uc_1427;
wire uc_1428;
wire uc_1429;
wire uc_1430;
wire uc_1431;
wire uc_1432;
wire uc_1433;
wire uc_1434;
wire uc_1435;
wire uc_1436;
wire uc_1437;
wire uc_1438;
wire uc_1439;
wire uc_1440;
wire uc_1441;
wire uc_1442;
wire uc_1443;
wire uc_1444;
wire uc_1445;
wire uc_1446;
wire uc_1447;
wire uc_1448;
wire uc_1449;
wire uc_1450;
wire uc_1451;
wire uc_1452;
wire uc_1453;
wire uc_1454;
wire uc_1455;
wire uc_1456;
wire uc_1457;
wire uc_1458;
wire uc_1459;
wire uc_1460;
wire uc_1461;
wire uc_1462;
wire uc_1463;
wire uc_1464;
wire uc_1465;
wire uc_1466;
wire uc_1467;
wire uc_1468;
wire uc_1469;
wire uc_1470;
wire uc_1471;
wire uc_1472;
wire uc_1473;
wire uc_1474;
wire uc_1475;
wire uc_1476;
wire uc_1477;
wire uc_1478;
wire uc_1479;
wire uc_1480;
wire uc_1481;
wire uc_1482;
wire uc_1483;
wire uc_1484;
wire uc_1485;
wire uc_1486;
wire uc_1487;
wire uc_1488;
wire uc_1489;
wire uc_1490;
wire uc_1491;
wire uc_1492;
wire uc_1493;
wire uc_1494;
wire uc_1495;
wire uc_1496;
wire uc_1497;
wire uc_1498;
wire uc_1499;
wire uc_1500;
wire uc_1501;
wire uc_1502;
wire uc_1503;
wire uc_1504;
wire uc_1505;
wire uc_1506;
wire uc_1507;
wire uc_1508;
wire uc_1509;
wire uc_1510;
wire uc_1511;
wire uc_1512;
wire uc_1513;
wire uc_1514;
wire uc_1515;
wire uc_1516;
wire uc_1517;
wire uc_1518;
wire uc_1519;
wire uc_1520;
wire uc_1521;
wire uc_1522;
wire uc_1523;
wire uc_1524;
wire uc_1525;
wire uc_1526;
wire uc_1527;
wire uc_1528;
wire uc_1529;
wire uc_1530;
wire uc_1531;
wire uc_1532;
wire uc_1533;
wire uc_1534;
wire uc_1535;
wire uc_1536;
wire uc_1537;
wire uc_1538;
wire uc_1539;
wire uc_1540;
wire uc_1541;
wire uc_1542;
wire uc_1543;
wire uc_1544;
wire uc_1545;
wire uc_1546;
wire uc_1547;
wire uc_1548;
wire uc_1549;
wire uc_1550;
wire uc_1551;
wire uc_1552;
wire uc_1553;
wire uc_1554;
wire uc_1555;
wire uc_1556;
wire uc_1557;
wire uc_1558;
wire uc_1559;
wire uc_1560;
wire uc_1561;
wire uc_1562;
wire uc_1563;
wire uc_1564;
wire uc_1565;
wire uc_1566;
wire uc_1567;
wire uc_1568;
wire uc_1569;
wire uc_1570;
wire uc_1571;
wire uc_1572;
wire uc_1573;
wire uc_1574;
wire uc_1575;
wire uc_1576;
wire uc_1577;
wire uc_1578;
wire uc_1579;
wire uc_1580;
wire uc_1581;
wire uc_1582;
wire uc_1583;
wire uc_1584;
wire uc_1585;
wire uc_1586;
wire uc_1587;
wire uc_1588;
wire uc_1589;
wire uc_1590;
wire uc_1591;
wire uc_1592;
wire uc_1593;
wire uc_1594;
wire uc_1595;
wire uc_1596;
wire uc_1597;
wire uc_1598;
wire uc_1599;
wire uc_1600;
wire uc_1601;
wire uc_1602;
wire uc_1603;
wire uc_1604;
wire uc_1605;
wire uc_1606;
wire uc_1607;
wire uc_1608;
wire uc_1609;
wire uc_1610;
wire uc_1611;
wire uc_1612;
wire uc_1613;
wire uc_1614;
wire uc_1615;
wire uc_1616;
wire uc_1617;
wire uc_1618;
wire uc_1619;
wire uc_1620;
wire uc_1621;
wire uc_1622;
wire uc_1623;
wire uc_1624;
wire uc_1625;
wire uc_1626;
wire uc_1627;
wire uc_1628;
wire uc_1629;
wire uc_1630;
wire uc_1631;
wire uc_1632;
wire uc_1633;
wire uc_1634;
wire uc_1635;
wire uc_1636;
wire uc_1637;
wire uc_1638;
wire uc_1639;
wire uc_1640;
wire uc_1641;
wire uc_1642;
wire uc_1643;
wire uc_1644;
wire uc_1645;
wire uc_1646;
wire uc_1647;
wire uc_1648;
wire uc_1649;
wire uc_1650;
wire uc_1651;
wire uc_1652;
wire uc_1653;
wire uc_1654;
wire uc_1655;
wire uc_1656;
wire uc_1657;
wire uc_1658;
wire uc_1659;
wire uc_1660;
wire uc_1661;
wire uc_1662;
wire uc_1663;
wire uc_1664;
wire uc_1665;
wire uc_1666;
wire uc_1667;
wire uc_1668;
wire uc_1669;
wire uc_1670;
wire uc_1671;
wire uc_1672;
wire uc_1673;
wire uc_1674;
wire uc_1675;
wire uc_1676;
wire uc_1677;
wire uc_1678;
wire uc_1679;
wire uc_1680;
wire uc_1681;
wire uc_1682;
wire uc_1683;
wire uc_1684;
wire uc_1685;
wire uc_1686;
wire uc_1687;
wire uc_1688;
wire uc_1689;
wire uc_1690;
wire uc_1691;
wire uc_1692;
wire uc_1693;
wire uc_1694;
wire uc_1695;
wire uc_1696;
wire uc_1697;
wire uc_1698;
wire uc_1699;
wire uc_1700;
wire uc_1701;
wire uc_1702;
wire uc_1703;
wire uc_1704;
wire uc_1705;
wire uc_1706;
wire uc_1707;
wire uc_1708;
wire uc_1709;
wire uc_1710;
wire uc_1711;
wire uc_1712;
wire uc_1713;
wire uc_1714;
wire uc_1715;
wire uc_1716;
wire uc_1717;
wire uc_1718;
wire uc_1719;
wire uc_1720;
wire uc_1721;
wire uc_1722;
wire uc_1723;
wire uc_1724;
wire uc_1725;
wire uc_1726;
wire uc_1727;
wire uc_1728;
wire uc_1729;
wire uc_1730;
wire uc_1731;
wire uc_1732;
wire uc_1733;
wire uc_1734;
wire uc_1735;
wire uc_1736;
wire uc_1737;
wire uc_1738;
wire uc_1739;
wire uc_1740;
wire uc_1741;
wire uc_1742;
wire uc_1743;
wire uc_1744;
wire uc_1745;
wire uc_1746;
wire uc_1747;
wire uc_1748;
wire uc_1749;
wire uc_1750;
wire uc_1751;
wire uc_1752;
wire uc_1753;
wire uc_1754;
wire uc_1755;
wire uc_1756;
wire uc_1757;
wire uc_1758;
wire uc_1759;
wire uc_1760;
wire uc_1761;
wire uc_1762;
wire uc_1763;
wire uc_1764;
wire uc_1765;
wire uc_1766;
wire uc_1767;
wire uc_1768;
wire uc_1769;
wire uc_1770;
wire uc_1771;
wire uc_1772;
wire uc_1773;
wire uc_1774;
wire uc_1775;
wire uc_1776;
wire uc_1777;
wire uc_1778;
wire uc_1779;
wire uc_1780;
wire uc_1781;
wire uc_1782;
wire uc_1783;
wire uc_1784;
wire uc_1785;
wire uc_1786;
wire uc_1787;
wire uc_1788;
wire uc_1789;
wire uc_1790;
wire uc_1791;
wire uc_1792;
wire uc_1793;
wire uc_1794;
wire uc_1795;
wire uc_1796;
wire uc_1797;
wire uc_1798;
wire uc_1799;
wire uc_1800;
wire uc_1801;
wire uc_1802;
wire uc_1803;
wire uc_1804;
wire uc_1805;
wire uc_1806;
wire uc_1807;
wire uc_1808;
wire uc_1809;
wire uc_1810;
wire uc_1811;
wire uc_1812;
wire uc_1813;
wire uc_1814;
wire uc_1815;
wire uc_1816;
wire uc_1817;
wire uc_1818;
wire uc_1819;
wire uc_1820;
wire uc_1821;
wire uc_1822;
wire uc_1823;
wire uc_1824;
wire uc_1825;
wire uc_1826;
wire uc_1827;
wire uc_1828;
wire uc_1829;
wire uc_1830;
wire uc_1831;
wire uc_1832;
wire uc_1833;
wire uc_1834;
wire uc_1835;
wire uc_1836;
wire uc_1837;
wire uc_1838;
wire uc_1839;
wire uc_1840;
wire uc_1841;
wire uc_1842;
wire uc_1843;
wire uc_1844;
wire uc_1845;
wire uc_1846;
wire uc_1847;
wire uc_1848;
wire uc_1849;
wire uc_1850;
wire uc_1851;
wire uc_1852;
wire uc_1853;
wire uc_1854;
wire uc_1855;
wire uc_1856;
wire uc_1857;
wire uc_1858;
wire uc_1859;
wire uc_1860;
wire uc_1861;
wire uc_1862;
wire uc_1863;
wire uc_1864;
wire uc_1865;
wire uc_1866;
wire uc_1867;
wire uc_1868;
wire uc_1869;
wire uc_1870;
wire uc_1871;
wire uc_1872;
wire uc_1873;
wire uc_1874;
wire uc_1875;
wire uc_1876;
wire uc_1877;
wire uc_1878;
wire uc_1879;
wire uc_1880;
wire uc_1881;
wire uc_1882;
wire uc_1883;
wire uc_1884;
wire uc_1885;
wire uc_1886;
wire uc_1887;
wire uc_1888;
wire uc_1889;
wire uc_1890;
wire uc_1891;
wire uc_1892;
wire uc_1893;
wire uc_1894;
wire uc_1895;
wire uc_1896;
wire uc_1897;
wire uc_1898;
wire uc_1899;
wire uc_1900;
wire uc_1901;
wire uc_1902;
wire uc_1903;
wire uc_1904;
wire uc_1905;
wire uc_1906;
wire uc_1907;
wire uc_1908;
wire uc_1909;
wire uc_1910;
wire uc_1911;
wire uc_1912;
wire uc_1913;
wire uc_1914;
wire uc_1915;
wire uc_1916;
wire uc_1917;
wire uc_1918;
wire uc_1919;
wire uc_1920;
wire uc_1921;
wire uc_1922;
wire uc_1923;
wire uc_1924;
wire uc_1925;
wire uc_1926;
wire uc_1927;
wire uc_1928;
wire uc_1929;
wire uc_1930;
wire uc_1931;
wire uc_1932;
wire uc_1933;
wire uc_1934;
wire uc_1935;
wire uc_1936;
wire uc_1937;
wire uc_1938;
wire uc_1939;
wire uc_1940;
wire uc_1941;
wire uc_1942;
wire uc_1943;
wire uc_1944;
wire uc_1945;
wire uc_1946;
wire uc_1947;
wire uc_1948;
wire uc_1949;
wire uc_1950;
wire uc_1951;
wire uc_1952;
wire uc_1953;
wire uc_1954;


WTM8 M1 (.Result ({\P[1][15] , \P[1][14] , \P[1][13] , \P[1][12] , \P[1][11] , \P[1][10] , 
    \P[1][9] , \P[1][8] , \P[1][7] , \P[1][6] , \P[1][5] , \P[1][4] , \P[1][3] , 
    \P[1][2] , \P[1][1] , \P[1][0] }), .A ({spw__n67, spw__n277, spw__n89, \a[4] , 
    \a[3] , \a[2] , \a[1] , A[0]}), .B ({\b[15] , \b[14] , spw__n226, \b[12] , \b[11] , 
    \b[10] , \b[9] , \b[8] }), .A_7_PP_0 (spw__n324), .A_5_PP_0 (spw__n90), .B_7_PP_0 (spw__n135)
    , .B_7_PP_1 (spw__n136), .B_7_PP_2 (spw__n139), .B_5_PP_0 (spw__n227), .B_5_PP_1 (spw__n228)
    , .B_5_PP_2 (spw__n229), .B_5_PP_3 (spw__n230), .A_7_PP_0PP_0 (spw__n325));
WTM8__2_1898 M8 (.Result ({\P[8][15] , \P[8][14] , \P[8][13] , \P[8][12] , \P[8][11] , 
    \P[8][10] , \P[8][9] , \P[8][8] , \Eight[1][23] , \Eight[1][22] , \Eight[1][21] , 
    \Eight[1][20] , \Eight[1][19] , \Eight[1][18] , \Eight[1][17] , \Eight[1][16] })
    , .A ({spw__n216, spw__n155, spw__n52, spw__n123, spw__n112, \a[18] , \a[17] , 
    \a[16] }), .B ({\b[7] , \b[6] , \b[5] , \b[4] , \b[3] , \b[2] , \b[1] , B[0]})
    , .A_5_PP_0 (spw__n53), .A_5_PP_1 (spw__n54), .A_4_PP_0 (spw__n124), .A_4_PP_1 (spw__n124)
    , .A_4_PP_2 (spw__n124), .A_4_PP_3 (spw__n124), .A_4_PP_4 (spw__n124), .B_5_PP_0 (spw__n314));
WTM8__2_1644 M9 (.Result ({\P[9][15] , \P[9][14] , \P[9][13] , \P[9][12] , \P[9][11] , 
    \P[9][10] , \P[9][9] , \P[9][8] , \P[9][7] , \P[9][6] , \P[9][5] , \P[9][4] , 
    \P[9][3] , \P[9][2] , \P[9][1] , \P[9][0] }), .A ({\a[23] , \a[22] , spw__n52, 
    spw__n123, spw__n112, \a[18] , \a[17] , \a[16] }), .B ({spw__n137, \b[14] , \b[13] , 
    \b[12] , \b[11] , \b[10] , \b[9] , \b[8] }), .A_4_PP_0 (spw__n123), .B_7_PP_0 (spw__n138)
    , .B_7_PP_1 (spw__n139), .A_6_PP_0 (spw__n152), .A_6_PP_1 (spw__n153), .A_6_PP_2 (spw__n154)
    , .A_6_PP_3 (spw__n155), .A_7_PP_0 (spw__n215), .A_7_PP_1 (spw__n216), .B_5_PP_0 (spw__n225));
adder64 A4 (.z ({uc_1908, uc_1909, uc_1910, uc_1911, uc_1912, uc_1913, uc_1914, uc_1915, 
    uc_1916, uc_1917, uc_1918, uc_1919, uc_1920, uc_1921, uc_1922, uc_1923, uc_1924, 
    uc_1925, uc_1926, uc_1927, uc_1928, uc_1929, uc_1930, \couple[4][40] , \couple[4][39] , 
    \couple[4][38] , \couple[4][37] , \couple[4][36] , \couple[4][35] , \couple[4][34] , 
    \couple[4][33] , \couple[4][32] , \couple[4][31] , \couple[4][30] , \couple[4][29] , 
    \couple[4][28] , \couple[4][27] , \couple[4][26] , \couple[4][25] , \couple[4][24] , 
    uc_1931, uc_1932, uc_1933, uc_1934, uc_1935, uc_1936, uc_1937, uc_1938, uc_1939, 
    uc_1940, uc_1941, uc_1942, uc_1943, uc_1944, uc_1945, uc_1946, uc_1947, uc_1948, 
    uc_1949, uc_1950, uc_1951, uc_1952, uc_1953, uc_1954}), .x ({uc_1804, uc_1805, 
    uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, uc_1811, uc_1812, uc_1813, uc_1814, 
    uc_1815, uc_1816, uc_1817, uc_1818, uc_1819, uc_1820, uc_1821, uc_1822, uc_1823, 
    uc_1824, uc_1825, uc_1826, uc_1827, uc_1828, uc_1829, uc_1830, uc_1831, uc_1832, 
    uc_1833, uc_1834, uc_1835, \P[8][15] , \P[8][14] , \P[8][13] , \P[8][12] , \P[8][11] , 
    \P[8][10] , \P[8][9] , \P[8][8] , uc_1836, uc_1837, uc_1838, uc_1839, uc_1840, 
    uc_1841, uc_1842, uc_1843, uc_1844, uc_1845, uc_1846, uc_1847, uc_1848, uc_1849, 
    uc_1850, uc_1851, uc_1852, uc_1853, uc_1854, uc_1855, uc_1856, uc_1857, uc_1858, 
    uc_1859}), .y ({uc_1860, uc_1861, uc_1862, uc_1863, uc_1864, uc_1865, uc_1866, 
    uc_1867, uc_1868, uc_1869, uc_1870, uc_1871, uc_1872, uc_1873, uc_1874, uc_1875, 
    uc_1876, uc_1877, uc_1878, uc_1879, uc_1880, uc_1881, uc_1882, uc_1883, \P[9][15] , 
    \P[9][14] , \P[9][13] , \P[9][12] , \P[9][11] , \P[9][10] , \P[9][9] , \P[9][8] , 
    \P[9][7] , \P[9][6] , \P[9][5] , \P[9][4] , \P[9][3] , \P[9][2] , \P[9][1] , 
    \P[9][0] , uc_1884, uc_1885, uc_1886, uc_1887, uc_1888, uc_1889, uc_1890, uc_1891, 
    uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, uc_1897, uc_1898, uc_1899, uc_1900, 
    uc_1901, uc_1902, uc_1903, uc_1904, uc_1905, uc_1906, uc_1907}));
WTM8__2_1390 M11 (.Result ({\P[11][15] , \P[11][14] , \P[11][13] , \P[11][12] , \P[11][11] , 
    \P[11][10] , \P[11][9] , \P[11][8] , \P[11][7] , \P[11][6] , \P[11][5] , \P[11][4] , 
    \P[11][3] , \P[11][2] , \P[11][1] , \P[11][0] }), .A ({\a[23] , \a[22] , \a[21] , 
    \a[20] , \a[19] , \a[18] , \a[17] , \a[16] }), .B ({\b[31] , \b[30] , \b[29] , 
    \b[28] , \b[27] , \b[26] , \b[25] , \b[24] }), .A_4_PP_0 (spw__n122));
adder64__2_3056 A5 (.z ({uc_1757, uc_1758, uc_1759, uc_1760, uc_1761, uc_1762, uc_1763, 
    \couple[5][56] , \couple[5][55] , \couple[5][54] , \couple[5][53] , \couple[5][52] , 
    \couple[5][51] , \couple[5][50] , \couple[5][49] , \couple[5][48] , \couple[5][47] , 
    \couple[5][46] , \couple[5][45] , \couple[5][44] , \couple[5][43] , \couple[5][42] , 
    \couple[5][41] , \couple[5][40] , uc_1764, uc_1765, uc_1766, uc_1767, uc_1768, 
    uc_1769, uc_1770, uc_1771, uc_1772, uc_1773, uc_1774, uc_1775, uc_1776, uc_1777, 
    uc_1778, uc_1779, uc_1780, uc_1781, uc_1782, uc_1783, uc_1784, uc_1785, uc_1786, 
    uc_1787, uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, uc_1793, uc_1794, uc_1795, 
    uc_1796, uc_1797, uc_1798, uc_1799, uc_1800, uc_1801, uc_1802, uc_1803}), .x ({
    uc_1653, uc_1654, uc_1655, uc_1656, uc_1657, uc_1658, uc_1659, uc_1660, uc_1661, 
    uc_1662, uc_1663, uc_1664, uc_1665, uc_1666, uc_1667, uc_1668, \P[10][15] , \P[10][14] , 
    \P[10][13] , \P[10][12] , \P[10][11] , \P[10][10] , \P[10][9] , \P[10][8] , uc_1669, 
    uc_1670, uc_1671, uc_1672, uc_1673, uc_1674, uc_1675, uc_1676, uc_1677, uc_1678, 
    uc_1679, uc_1680, uc_1681, uc_1682, uc_1683, uc_1684, uc_1685, uc_1686, uc_1687, 
    uc_1688, uc_1689, uc_1690, uc_1691, uc_1692, uc_1693, uc_1694, uc_1695, uc_1696, 
    uc_1697, uc_1698, uc_1699, uc_1700, uc_1701, uc_1702, uc_1703, uc_1704, uc_1705, 
    uc_1706, uc_1707, uc_1708}), .y ({uc_1709, uc_1710, uc_1711, uc_1712, uc_1713, 
    uc_1714, uc_1715, uc_1716, \P[11][15] , \P[11][14] , \P[11][13] , \P[11][12] , 
    \P[11][11] , \P[11][10] , \P[11][9] , \P[11][8] , \P[11][7] , \P[11][6] , \P[11][5] , 
    \P[11][4] , \P[11][3] , \P[11][2] , \P[11][1] , \P[11][0] , uc_1717, uc_1718, 
    uc_1719, uc_1720, uc_1721, uc_1722, uc_1723, uc_1724, uc_1725, uc_1726, uc_1727, 
    uc_1728, uc_1729, uc_1730, uc_1731, uc_1732, uc_1733, uc_1734, uc_1735, uc_1736, 
    uc_1737, uc_1738, uc_1739, uc_1740, uc_1741, uc_1742, uc_1743, uc_1744, uc_1745, 
    uc_1746, uc_1747, uc_1748, uc_1749, uc_1750, uc_1751, uc_1752, uc_1753, uc_1754, 
    uc_1755, uc_1756}));
adder64__2_2863 A10 (.z ({uc_1615, uc_1616, uc_1617, uc_1618, uc_1619, uc_1620, \Quadruple[2][57] , 
    \Quadruple[2][56] , \Quadruple[2][55] , \Quadruple[2][54] , \Quadruple[2][53] , 
    \Quadruple[2][52] , \Quadruple[2][51] , \Quadruple[2][50] , \Quadruple[2][49] , 
    \Quadruple[2][48] , \Quadruple[2][47] , \Quadruple[2][46] , \Quadruple[2][45] , 
    \Quadruple[2][44] , \Quadruple[2][43] , \Quadruple[2][42] , \Quadruple[2][41] , 
    \Quadruple[2][40] , \Quadruple[2][39] , \Quadruple[2][38] , \Quadruple[2][37] , 
    \Quadruple[2][36] , \Quadruple[2][35] , \Quadruple[2][34] , \Quadruple[2][33] , 
    \Quadruple[2][32] , uc_1621, uc_1622, uc_1623, uc_1624, uc_1625, uc_1626, uc_1627, 
    uc_1628, uc_1629, uc_1630, uc_1631, uc_1632, uc_1633, uc_1634, uc_1635, uc_1636, 
    uc_1637, uc_1638, uc_1639, uc_1640, uc_1641, uc_1642, uc_1643, uc_1644, uc_1645, 
    uc_1646, uc_1647, uc_1648, uc_1649, uc_1650, uc_1651, uc_1652}), .x ({uc_1521, 
    uc_1522, uc_1523, uc_1524, uc_1525, uc_1526, uc_1527, uc_1528, uc_1529, uc_1530, 
    uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, uc_1538, uc_1539, 
    uc_1540, uc_1541, uc_1542, uc_1543, \couple[4][40] , \couple[4][39] , \couple[4][38] , 
    \couple[4][37] , \couple[4][36] , \couple[4][35] , \couple[4][34] , \couple[4][33] , 
    \couple[4][32] , uc_1544, uc_1545, uc_1546, uc_1547, uc_1548, uc_1549, uc_1550, 
    uc_1551, uc_1552, uc_1553, uc_1554, uc_1555, uc_1556, uc_1557, uc_1558, uc_1559, 
    uc_1560, uc_1561, uc_1562, uc_1563, uc_1564, uc_1565, uc_1566, uc_1567, uc_1568, 
    uc_1569, uc_1570, uc_1571, uc_1572, uc_1573, uc_1574, uc_1575}), .y ({uc_1576, 
    uc_1577, uc_1578, uc_1579, uc_1580, uc_1581, uc_1582, \couple[5][56] , \couple[5][55] , 
    \couple[5][54] , \couple[5][53] , \couple[5][52] , \couple[5][51] , \couple[5][50] , 
    \couple[5][49] , \couple[5][48] , \couple[5][47] , \couple[5][46] , \couple[5][45] , 
    \couple[5][44] , \couple[5][43] , \couple[5][42] , \couple[5][41] , \couple[5][40] , 
    \P[10][7] , \P[10][6] , \P[10][5] , \P[10][4] , \P[10][3] , \P[10][2] , \P[10][1] , 
    \P[10][0] , uc_1583, uc_1584, uc_1585, uc_1586, uc_1587, uc_1588, uc_1589, uc_1590, 
    uc_1591, uc_1592, uc_1593, uc_1594, uc_1595, uc_1596, uc_1597, uc_1598, uc_1599, 
    uc_1600, uc_1601, uc_1602, uc_1603, uc_1604, uc_1605, uc_1606, uc_1607, uc_1608, 
    uc_1609, uc_1610, uc_1611, uc_1612, uc_1613, uc_1614}));
WTM8__2_1136 M12 (.Result ({\P[12][15] , \P[12][14] , \P[12][13] , \P[12][12] , \P[12][11] , 
    \P[12][10] , \P[12][9] , \P[12][8] , \P[12][7] , \P[12][6] , \P[12][5] , \P[12][4] , 
    \P[12][3] , \P[12][2] , \P[12][1] , \P[12][0] }), .A ({\a[31] , \a[30] , \a[29] , 
    \a[28] , \a[27] , \a[26] , \a[25] , \a[24] }), .B ({\b[7] , \b[6] , spw__n314, 
    \b[4] , \b[3] , \b[2] , \b[1] , B[0]}));
adder64__2_2670 A13 (.z ({\Eight[1][63] , \Eight[1][62] , \Eight[1][61] , \Eight[1][60] , 
    \Eight[1][59] , \Eight[1][58] , \Eight[1][57] , \Eight[1][56] , \Eight[1][55] , 
    \Eight[1][54] , \Eight[1][53] , \Eight[1][52] , \Eight[1][51] , \Eight[1][50] , 
    \Eight[1][49] , \Eight[1][48] , \Eight[1][47] , \Eight[1][46] , \Eight[1][45] , 
    \Eight[1][44] , \Eight[1][43] , \Eight[1][42] , \Eight[1][41] , \Eight[1][40] , 
    \Eight[1][39] , \Eight[1][38] , \Eight[1][37] , \Eight[1][36] , \Eight[1][35] , 
    \Eight[1][34] , \Eight[1][33] , \Eight[1][32] , \Eight[1][31] , \Eight[1][30] , 
    \Eight[1][29] , \Eight[1][28] , \Eight[1][27] , \Eight[1][26] , \Eight[1][25] , 
    \Eight[1][24] , uc_1497, uc_1498, uc_1499, uc_1500, uc_1501, uc_1502, uc_1503, 
    uc_1504, uc_1505, uc_1506, uc_1507, uc_1508, uc_1509, uc_1510, uc_1511, uc_1512, 
    uc_1513, uc_1514, uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, uc_1520}), .x ({
    uc_1443, uc_1444, uc_1445, uc_1446, uc_1447, uc_1448, \Quadruple[2][57] , \Quadruple[2][56] , 
    \Quadruple[2][55] , \Quadruple[2][54] , \Quadruple[2][53] , \Quadruple[2][52] , 
    \Quadruple[2][51] , \Quadruple[2][50] , \Quadruple[2][49] , \Quadruple[2][48] , 
    \Quadruple[2][47] , \Quadruple[2][46] , \Quadruple[2][45] , \Quadruple[2][44] , 
    \Quadruple[2][43] , \Quadruple[2][42] , \Quadruple[2][41] , \Quadruple[2][40] , 
    \Quadruple[2][39] , \Quadruple[2][38] , \Quadruple[2][37] , \Quadruple[2][36] , 
    \Quadruple[2][35] , \Quadruple[2][34] , \Quadruple[2][33] , \Quadruple[2][32] , 
    \couple[4][31] , \couple[4][30] , \couple[4][29] , \couple[4][28] , \couple[4][27] , 
    \couple[4][26] , \couple[4][25] , \couple[4][24] , uc_1449, uc_1450, uc_1451, 
    uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, uc_1458, uc_1459, uc_1460, 
    uc_1461, uc_1462, uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, 
    uc_1470, uc_1471, uc_1472}), .y ({\Quadruple[3][63] , \Quadruple[3][62] , \Quadruple[3][61] , 
    \Quadruple[3][60] , \Quadruple[3][59] , \Quadruple[3][58] , \Quadruple[3][57] , 
    \Quadruple[3][56] , \Quadruple[3][55] , \Quadruple[3][54] , \Quadruple[3][53] , 
    \Quadruple[3][52] , \Quadruple[3][51] , \Quadruple[3][50] , \Quadruple[3][49] , 
    \Quadruple[3][48] , \Quadruple[3][47] , \Quadruple[3][46] , \Quadruple[3][45] , 
    \Quadruple[3][44] , \Quadruple[3][43] , \Quadruple[3][42] , \Quadruple[3][41] , 
    \Quadruple[3][40] , \couple[6][39] , \couple[6][38] , \couple[6][37] , \couple[6][36] , 
    \couple[6][35] , \couple[6][34] , \couple[6][33] , \couple[6][32] , \P[12][7] , 
    \P[12][6] , \P[12][5] , \P[12][4] , \P[12][3] , \P[12][2] , \P[12][1] , \P[12][0] , 
    uc_1473, uc_1474, uc_1475, uc_1476, uc_1477, uc_1478, uc_1479, uc_1480, uc_1481, 
    uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, uc_1488, uc_1489, uc_1490, 
    uc_1491, uc_1492, uc_1493, uc_1494, uc_1495, uc_1496}));
adder64__2_2477 A11 (.z ({\Quadruple[3][63] , \Quadruple[3][62] , \Quadruple[3][61] , 
    \Quadruple[3][60] , \Quadruple[3][59] , \Quadruple[3][58] , \Quadruple[3][57] , 
    \Quadruple[3][56] , \Quadruple[3][55] , \Quadruple[3][54] , \Quadruple[3][53] , 
    \Quadruple[3][52] , \Quadruple[3][51] , \Quadruple[3][50] , \Quadruple[3][49] , 
    \Quadruple[3][48] , \Quadruple[3][47] , \Quadruple[3][46] , \Quadruple[3][45] , 
    \Quadruple[3][44] , \Quadruple[3][43] , \Quadruple[3][42] , \Quadruple[3][41] , 
    \Quadruple[3][40] , uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, uc_1408, uc_1409, 
    uc_1410, uc_1411, uc_1412, uc_1413, uc_1414, uc_1415, uc_1416, uc_1417, uc_1418, 
    uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, uc_1427, 
    uc_1428, uc_1429, uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, uc_1435, uc_1436, 
    uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442}), .x ({uc_1308, uc_1309, 
    uc_1310, uc_1311, uc_1312, uc_1313, uc_1314, uc_1315, uc_1316, uc_1317, uc_1318, 
    uc_1319, uc_1320, uc_1321, uc_1322, \couple[6][48] , \couple[6][47] , \couple[6][46] , 
    \couple[6][45] , \couple[6][44] , \couple[6][43] , \couple[6][42] , \couple[6][41] , 
    \couple[6][40] , uc_1323, uc_1324, uc_1325, uc_1326, uc_1327, uc_1328, uc_1329, 
    uc_1330, uc_1331, uc_1332, uc_1333, uc_1334, uc_1335, uc_1336, uc_1337, uc_1338, 
    uc_1339, uc_1340, uc_1341, uc_1342, uc_1343, uc_1344, uc_1345, uc_1346, uc_1347, 
    uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, uc_1353, uc_1354, uc_1355, uc_1356, 
    uc_1357, uc_1358, uc_1359, uc_1360, uc_1361, uc_1362}), .y ({\couple[7][63] , 
    \couple[7][62] , \couple[7][61] , \couple[7][60] , \couple[7][59] , \couple[7][58] , 
    \couple[7][57] , \couple[7][56] , \couple[7][55] , \couple[7][54] , \couple[7][53] , 
    \couple[7][52] , \couple[7][51] , \couple[7][50] , \couple[7][49] , \couple[7][48] , 
    \P[14][7] , \P[14][6] , \P[14][5] , \P[14][4] , \P[14][3] , \P[14][2] , \P[14][1] , 
    \P[14][0] , uc_1363, uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, 
    uc_1371, uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, uc_1378, uc_1379, 
    uc_1380, uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, 
    uc_1389, uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396, uc_1397, 
    uc_1398, uc_1399, uc_1400, uc_1401, uc_1402}));
adder64__2_2284 A7 (.z ({\couple[7][63] , \couple[7][62] , \couple[7][61] , \couple[7][60] , 
    \couple[7][59] , \couple[7][58] , \couple[7][57] , \couple[7][56] , \couple[7][55] , 
    \couple[7][54] , \couple[7][53] , \couple[7][52] , \couple[7][51] , \couple[7][50] , 
    \couple[7][49] , \couple[7][48] , uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, 
    uc_1265, uc_1266, uc_1267, uc_1268, uc_1269, uc_1270, uc_1271, uc_1272, uc_1273, 
    uc_1274, uc_1275, uc_1276, uc_1277, uc_1278, uc_1279, uc_1280, uc_1281, uc_1282, 
    uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, uc_1288, uc_1289, uc_1290, uc_1291, 
    uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, 
    uc_1301, uc_1302, uc_1303, uc_1304, uc_1305, uc_1306, uc_1307}), .x ({uc_1156, 
    uc_1157, uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, \P[14][15] , \P[14][14] , 
    \P[14][13] , \P[14][12] , \P[14][11] , \P[14][10] , \P[14][9] , \P[14][8] , uc_1164, 
    uc_1165, uc_1166, uc_1167, uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, 
    uc_1174, uc_1175, uc_1176, uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, 
    uc_1183, uc_1184, uc_1185, uc_1186, uc_1187, uc_1188, uc_1189, uc_1190, uc_1191, 
    uc_1192, uc_1193, uc_1194, uc_1195, uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, 
    uc_1201, uc_1202, uc_1203, uc_1204, uc_1205, uc_1206, uc_1207, uc_1208, uc_1209, 
    uc_1210, uc_1211}), .y ({\P[15][15] , \P[15][14] , \P[15][13] , \P[15][12] , 
    \P[15][11] , \P[15][10] , \P[15][9] , \P[15][8] , \P[15][7] , \P[15][6] , \P[15][5] , 
    \P[15][4] , \P[15][3] , \P[15][2] , \P[15][1] , \P[15][0] , uc_1212, uc_1213, 
    uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, 
    uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, 
    uc_1232, uc_1233, uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, uc_1239, uc_1240, 
    uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, uc_1249, 
    uc_1250, uc_1251, uc_1252, uc_1253, uc_1254, uc_1255, uc_1256, uc_1257, uc_1258, 
    uc_1259}));
WTM8__2_882 M15 (.Result ({\P[15][15] , \P[15][14] , \P[15][13] , \P[15][12] , \P[15][11] , 
    \P[15][10] , \P[15][9] , \P[15][8] , \P[15][7] , \P[15][6] , \P[15][5] , \P[15][4] , 
    \P[15][3] , \P[15][2] , \P[15][1] , \P[15][0] }), .A ({\a[31] , \a[30] , \a[29] , 
    \a[28] , \a[27] , \a[26] , \a[25] , \a[24] }), .B ({\b[31] , \b[30] , \b[29] , 
    \b[28] , \b[27] , \b[26] , \b[25] , \b[24] }));
WTM8__2_628 M13 (.Result ({\P[13][15] , \P[13][14] , \P[13][13] , \P[13][12] , \P[13][11] , 
    \P[13][10] , \P[13][9] , \P[13][8] , \P[13][7] , \P[13][6] , \P[13][5] , \P[13][4] , 
    \P[13][3] , \P[13][2] , \P[13][1] , \P[13][0] }), .A ({\a[31] , \a[30] , \a[29] , 
    \a[28] , \a[27] , \a[26] , \a[25] , \a[24] }), .B ({spw__n137, \b[14] , \b[13] , 
    \b[12] , \b[11] , \b[10] , \b[9] , \b[8] }));
adder64__2_2091 A6 (.z ({uc_1109, uc_1110, uc_1111, uc_1112, uc_1113, uc_1114, uc_1115, 
    uc_1116, uc_1117, uc_1118, uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, \couple[6][48] , 
    \couple[6][47] , \couple[6][46] , \couple[6][45] , \couple[6][44] , \couple[6][43] , 
    \couple[6][42] , \couple[6][41] , \couple[6][40] , \couple[6][39] , \couple[6][38] , 
    \couple[6][37] , \couple[6][36] , \couple[6][35] , \couple[6][34] , \couple[6][33] , 
    \couple[6][32] , uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, 
    uc_1131, uc_1132, uc_1133, uc_1134, uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, 
    uc_1140, uc_1141, uc_1142, uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, uc_1148, 
    uc_1149, uc_1150, uc_1151, uc_1152, uc_1153, uc_1154, uc_1155}), .x ({uc_1005, 
    uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, uc_1013, uc_1014, 
    uc_1015, uc_1016, uc_1017, uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, 
    uc_1024, uc_1025, uc_1026, uc_1027, uc_1028, \P[12][15] , \P[12][14] , \P[12][13] , 
    \P[12][12] , \P[12][11] , \P[12][10] , \P[12][9] , \P[12][8] , uc_1029, uc_1030, 
    uc_1031, uc_1032, uc_1033, uc_1034, uc_1035, uc_1036, uc_1037, uc_1038, uc_1039, 
    uc_1040, uc_1041, uc_1042, uc_1043, uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, 
    uc_1049, uc_1050, uc_1051, uc_1052, uc_1053, uc_1054, uc_1055, uc_1056, uc_1057, 
    uc_1058, uc_1059, uc_1060}), .y ({uc_1061, uc_1062, uc_1063, uc_1064, uc_1065, 
    uc_1066, uc_1067, uc_1068, uc_1069, uc_1070, uc_1071, uc_1072, uc_1073, uc_1074, 
    uc_1075, uc_1076, \P[13][15] , \P[13][14] , \P[13][13] , \P[13][12] , \P[13][11] , 
    \P[13][10] , \P[13][9] , \P[13][8] , \P[13][7] , \P[13][6] , \P[13][5] , \P[13][4] , 
    \P[13][3] , \P[13][2] , \P[13][1] , \P[13][0] , uc_1077, uc_1078, uc_1079, uc_1080, 
    uc_1081, uc_1082, uc_1083, uc_1084, uc_1085, uc_1086, uc_1087, uc_1088, uc_1089, 
    uc_1090, uc_1091, uc_1092, uc_1093, uc_1094, uc_1095, uc_1096, uc_1097, uc_1098, 
    uc_1099, uc_1100, uc_1101, uc_1102, uc_1103, uc_1104, uc_1105, uc_1106, uc_1107, 
    uc_1108}));
MUX2_X2 i_0_0_125 (.Z (Result[63]), .A (n_0_62), .B (\out[63] ), .S (sps__n1));
MUX2_X1 i_0_0_124 (.Z (Result[62]), .A (n_0_124), .B (\out[62] ), .S (sps__n1));
MUX2_X2 i_0_0_123 (.Z (Result[61]), .A (n_0_123), .B (\out[61] ), .S (sps__n1));
MUX2_X1 i_0_0_122 (.Z (Result[60]), .A (n_0_122), .B (\out[60] ), .S (sps__n1));
MUX2_X1 i_0_0_121 (.Z (Result[59]), .A (n_0_121), .B (\out[59] ), .S (sps__n1));
MUX2_X1 i_0_0_120 (.Z (Result[58]), .A (n_0_120), .B (\out[58] ), .S (sps__n1));
MUX2_X1 i_0_0_119 (.Z (Result[57]), .A (n_0_119), .B (\out[57] ), .S (sps__n1));
MUX2_X1 i_0_0_118 (.Z (Result[56]), .A (n_0_118), .B (\out[56] ), .S (sps__n1));
MUX2_X1 i_0_0_117 (.Z (Result[55]), .A (n_0_117), .B (\out[55] ), .S (sps__n1));
MUX2_X1 i_0_0_116 (.Z (Result[54]), .A (n_0_116), .B (\out[54] ), .S (sps__n1));
MUX2_X1 i_0_0_115 (.Z (Result[53]), .A (n_0_115), .B (\out[53] ), .S (sps__n1));
MUX2_X1 i_0_0_114 (.Z (Result[52]), .A (n_0_114), .B (\out[52] ), .S (sps__n1));
MUX2_X1 i_0_0_113 (.Z (Result[51]), .A (n_0_113), .B (\out[51] ), .S (sps__n1));
MUX2_X1 i_0_0_112 (.Z (Result[50]), .A (n_0_112), .B (\out[50] ), .S (sps__n1));
MUX2_X1 i_0_0_111 (.Z (Result[49]), .A (n_0_111), .B (\out[49] ), .S (sps__n1));
MUX2_X1 i_0_0_110 (.Z (Result[48]), .A (n_0_110), .B (\out[48] ), .S (sps__n1));
MUX2_X1 i_0_0_109 (.Z (Result[47]), .A (n_0_109), .B (\out[47] ), .S (sps__n1));
MUX2_X1 i_0_0_108 (.Z (Result[46]), .A (n_0_108), .B (\out[46] ), .S (sps__n1));
MUX2_X1 i_0_0_107 (.Z (Result[45]), .A (n_0_107), .B (\out[45] ), .S (sps__n1));
MUX2_X1 i_0_0_106 (.Z (Result[44]), .A (n_0_106), .B (\out[44] ), .S (sps__n1));
MUX2_X1 i_0_0_105 (.Z (Result[43]), .A (n_0_105), .B (\out[43] ), .S (sps__n1));
MUX2_X1 i_0_0_104 (.Z (Result[42]), .A (n_0_104), .B (\out[42] ), .S (sps__n1));
MUX2_X1 i_0_0_103 (.Z (Result[41]), .A (n_0_103), .B (\out[41] ), .S (sps__n1));
MUX2_X1 i_0_0_102 (.Z (Result[40]), .A (n_0_102), .B (\out[40] ), .S (sps__n1));
MUX2_X1 i_0_0_101 (.Z (Result[39]), .A (n_0_101), .B (\out[39] ), .S (sps__n1));
MUX2_X1 i_0_0_100 (.Z (Result[38]), .A (n_0_100), .B (\out[38] ), .S (sps__n1));
MUX2_X1 i_0_0_99 (.Z (Result[37]), .A (n_0_99), .B (\out[37] ), .S (sps__n1));
MUX2_X1 i_0_0_98 (.Z (Result[36]), .A (n_0_98), .B (\out[36] ), .S (sps__n1));
MUX2_X1 i_0_0_97 (.Z (Result[35]), .A (n_0_97), .B (\out[35] ), .S (sps__n1));
MUX2_X1 i_0_0_96 (.Z (Result[34]), .A (n_0_96), .B (\out[34] ), .S (sps__n1));
MUX2_X1 i_0_0_95 (.Z (Result[33]), .A (n_0_95), .B (\out[33] ), .S (sps__n1));
MUX2_X1 i_0_0_94 (.Z (Result[32]), .A (n_0_94), .B (\out[32] ), .S (sps__n1));
MUX2_X1 i_0_0_93 (.Z (Result[31]), .A (n_0_93), .B (\out[31] ), .S (sps__n1));
MUX2_X1 i_0_0_92 (.Z (Result[30]), .A (n_0_92), .B (\out[30] ), .S (sps__n1));
MUX2_X1 i_0_0_91 (.Z (Result[29]), .A (n_0_91), .B (\out[29] ), .S (sps__n1));
MUX2_X1 i_0_0_90 (.Z (Result[28]), .A (n_0_90), .B (\out[28] ), .S (sps__n1));
MUX2_X1 i_0_0_89 (.Z (Result[27]), .A (n_0_89), .B (\out[27] ), .S (sps__n1));
MUX2_X1 i_0_0_88 (.Z (Result[26]), .A (n_0_88), .B (\out[26] ), .S (sps__n1));
MUX2_X1 i_0_0_87 (.Z (Result[25]), .A (n_0_87), .B (\out[25] ), .S (sps__n1));
MUX2_X1 i_0_0_86 (.Z (Result[24]), .A (n_0_86), .B (\out[24] ), .S (sps__n1));
MUX2_X1 i_0_0_85 (.Z (Result[23]), .A (n_0_85), .B (\out[23] ), .S (sps__n1));
MUX2_X1 i_0_0_84 (.Z (Result[22]), .A (n_0_84), .B (\out[22] ), .S (sps__n1));
MUX2_X1 i_0_0_83 (.Z (Result[21]), .A (n_0_83), .B (\out[21] ), .S (sps__n1));
MUX2_X1 i_0_0_82 (.Z (Result[20]), .A (n_0_82), .B (\out[20] ), .S (sps__n1));
MUX2_X1 i_0_0_81 (.Z (Result[19]), .A (n_0_81), .B (\out[19] ), .S (sps__n1));
MUX2_X1 i_0_0_80 (.Z (Result[18]), .A (n_0_80), .B (\out[18] ), .S (sps__n1));
MUX2_X1 i_0_0_79 (.Z (Result[17]), .A (n_0_79), .B (\out[17] ), .S (sps__n1));
MUX2_X1 i_0_0_78 (.Z (Result[16]), .A (n_0_78), .B (\out[16] ), .S (sps__n1));
MUX2_X1 i_0_0_77 (.Z (Result[15]), .A (n_0_77), .B (\Eight[0][15] ), .S (sps__n1));
MUX2_X1 i_0_0_76 (.Z (Result[14]), .A (n_0_76), .B (\Eight[0][14] ), .S (sps__n1));
MUX2_X1 i_0_0_75 (.Z (Result[13]), .A (n_0_75), .B (\Eight[0][13] ), .S (sps__n1));
MUX2_X1 i_0_0_74 (.Z (Result[12]), .A (n_0_74), .B (\Eight[0][12] ), .S (sps__n1));
MUX2_X1 i_0_0_73 (.Z (Result[11]), .A (n_0_73), .B (\Eight[0][11] ), .S (sps__n1));
MUX2_X1 i_0_0_72 (.Z (Result[10]), .A (n_0_72), .B (\Eight[0][10] ), .S (sps__n1));
MUX2_X1 i_0_0_71 (.Z (Result[9]), .A (n_0_71), .B (\Eight[0][9] ), .S (sps__n1));
MUX2_X1 i_0_0_70 (.Z (Result[8]), .A (n_0_70), .B (\Eight[0][8] ), .S (sps__n1));
MUX2_X1 i_0_0_69 (.Z (Result[7]), .A (n_0_69), .B (\P[0][7] ), .S (sps__n1));
MUX2_X1 i_0_0_68 (.Z (Result[6]), .A (n_0_68), .B (\P[0][6] ), .S (sps__n1));
MUX2_X1 i_0_0_67 (.Z (Result[5]), .A (n_0_67), .B (\P[0][5] ), .S (sps__n1));
MUX2_X1 i_0_0_66 (.Z (Result[4]), .A (n_0_66), .B (\P[0][4] ), .S (sps__n1));
MUX2_X1 i_0_0_65 (.Z (Result[3]), .A (n_0_65), .B (\P[0][3] ), .S (sps__n1));
MUX2_X1 i_0_0_64 (.Z (Result[2]), .A (n_0_64), .B (\P[0][2] ), .S (sps__n1));
MUX2_X1 i_0_0_63 (.Z (Result[1]), .A (n_0_63), .B (\P[0][1] ), .S (sps__n1));
XNOR2_X1 i_0_0_62 (.ZN (n_0_0_0), .A (B[31]), .B (A[31]));
AND2_X2 i_0_0_61 (.ZN (\a[31] ), .A1 (n_0_61), .A2 (A[31]));
MUX2_X2 i_0_0_60 (.Z (\a[30] ), .A (A[30]), .B (n_0_60), .S (A[31]));
MUX2_X2 i_0_0_59 (.Z (\a[29] ), .A (A[29]), .B (n_0_59), .S (A[31]));
MUX2_X2 i_0_0_58 (.Z (\a[28] ), .A (A[28]), .B (n_0_58), .S (A[31]));
MUX2_X2 i_0_0_57 (.Z (\a[27] ), .A (A[27]), .B (n_0_57), .S (A[31]));
MUX2_X2 i_0_0_56 (.Z (\a[26] ), .A (A[26]), .B (n_0_56), .S (A[31]));
MUX2_X1 i_0_0_55 (.Z (\a[25] ), .A (A[25]), .B (n_0_55), .S (A[31]));
MUX2_X1 i_0_0_54 (.Z (\a[24] ), .A (A[24]), .B (n_0_54), .S (A[31]));
MUX2_X2 i_0_0_53 (.Z (spw__n216), .A (A[23]), .B (n_0_53), .S (A[31]));
MUX2_X2 i_0_0_52 (.Z (spw__n155), .A (A[22]), .B (n_0_52), .S (A[31]));
MUX2_X1 i_0_0_51 (.Z (spw__n54), .A (A[21]), .B (n_0_51), .S (A[31]));
MUX2_X1 i_0_0_50 (.Z (spw__n124), .A (A[20]), .B (n_0_50), .S (A[31]));
MUX2_X1 i_0_0_49 (.Z (spw__n113), .A (A[19]), .B (n_0_49), .S (A[31]));
MUX2_X2 i_0_0_48 (.Z (spw__n384), .A (A[18]), .B (n_0_48), .S (A[31]));
MUX2_X2 i_0_0_47 (.Z (\a[17] ), .A (A[17]), .B (n_0_47), .S (A[31]));
MUX2_X2 i_0_0_46 (.Z (\a[16] ), .A (A[16]), .B (n_0_46), .S (A[31]));
MUX2_X1 i_0_0_45 (.Z (spw__n184), .A (A[15]), .B (n_0_45), .S (A[31]));
MUX2_X1 i_0_0_44 (.Z (spw__n167), .A (A[14]), .B (n_0_44), .S (A[31]));
MUX2_X1 i_0_0_43 (.Z (spw__n81), .A (A[13]), .B (n_0_43), .S (A[31]));
MUX2_X2 i_0_0_42 (.Z (\a[12] ), .A (A[12]), .B (n_0_42), .S (A[31]));
MUX2_X2 i_0_0_41 (.Z (\a[11] ), .A (A[11]), .B (n_0_41), .S (A[31]));
MUX2_X2 i_0_0_40 (.Z (\a[10] ), .A (A[10]), .B (n_0_40), .S (A[31]));
MUX2_X2 i_0_0_39 (.Z (\a[9] ), .A (A[9]), .B (n_0_39), .S (A[31]));
MUX2_X2 i_0_0_38 (.Z (\a[8] ), .A (A[8]), .B (n_0_38), .S (A[31]));
MUX2_X2 i_0_0_37 (.Z (spw__n325), .A (A[7]), .B (n_0_37), .S (A[31]));
MUX2_X2 i_0_0_36 (.Z (spw__n278), .A (A[6]), .B (n_0_36), .S (A[31]));
MUX2_X2 i_0_0_35 (.Z (spt__n12), .A (A[5]), .B (n_0_35), .S (A[31]));
MUX2_X2 i_0_0_34 (.Z (\a[4] ), .A (A[4]), .B (n_0_34), .S (A[31]));
MUX2_X2 i_0_0_33 (.Z (\a[3] ), .A (A[3]), .B (n_0_33), .S (A[31]));
MUX2_X2 i_0_0_32 (.Z (\a[2] ), .A (A[2]), .B (n_0_32), .S (A[31]));
MUX2_X1 i_0_0_31 (.Z (\a[1] ), .A (A[1]), .B (n_0_31), .S (A[31]));
AND2_X1 i_0_0_30 (.ZN (\b[31] ), .A1 (n_0_30), .A2 (B[31]));
MUX2_X1 i_0_0_29 (.Z (\b[30] ), .A (B[30]), .B (n_0_29), .S (B[31]));
MUX2_X2 i_0_0_28 (.Z (\b[29] ), .A (B[29]), .B (n_0_28), .S (B[31]));
MUX2_X1 i_0_0_27 (.Z (\b[28] ), .A (B[28]), .B (n_0_27), .S (B[31]));
MUX2_X1 i_0_0_26 (.Z (\b[27] ), .A (B[27]), .B (n_0_26), .S (B[31]));
MUX2_X1 i_0_0_25 (.Z (\b[26] ), .A (B[26]), .B (n_0_25), .S (B[31]));
MUX2_X1 i_0_0_24 (.Z (\b[25] ), .A (B[25]), .B (n_0_24), .S (B[31]));
MUX2_X1 i_0_0_23 (.Z (\b[24] ), .A (B[24]), .B (n_0_23), .S (B[31]));
MUX2_X2 i_0_0_22 (.Z (\b[23] ), .A (B[23]), .B (n_0_22), .S (B[31]));
MUX2_X2 i_0_0_21 (.Z (\b[22] ), .A (B[22]), .B (n_0_21), .S (B[31]));
MUX2_X2 i_0_0_20 (.Z (\b[21] ), .A (B[21]), .B (n_0_20), .S (B[31]));
MUX2_X2 i_0_0_19 (.Z (\b[20] ), .A (B[20]), .B (n_0_19), .S (B[31]));
MUX2_X2 i_0_0_18 (.Z (\b[19] ), .A (B[19]), .B (n_0_18), .S (B[31]));
MUX2_X2 i_0_0_17 (.Z (\b[18] ), .A (B[18]), .B (n_0_17), .S (B[31]));
MUX2_X1 i_0_0_16 (.Z (\b[17] ), .A (B[17]), .B (n_0_16), .S (B[31]));
MUX2_X1 i_0_0_15 (.Z (\b[16] ), .A (B[16]), .B (n_0_15), .S (B[31]));
MUX2_X1 i_0_0_14 (.Z (spw__n139), .A (B[15]), .B (n_0_14), .S (B[31]));
MUX2_X2 i_0_0_13 (.Z (\b[14] ), .A (B[14]), .B (n_0_13), .S (B[31]));
MUX2_X2 i_0_0_12 (.Z (spw__n230), .A (B[13]), .B (n_0_12), .S (B[31]));
MUX2_X2 i_0_0_11 (.Z (\b[12] ), .A (B[12]), .B (n_0_11), .S (B[31]));
MUX2_X2 i_0_0_10 (.Z (\b[11] ), .A (B[11]), .B (n_0_10), .S (B[31]));
MUX2_X2 i_0_0_9 (.Z (\b[10] ), .A (B[10]), .B (n_0_9), .S (B[31]));
MUX2_X2 i_0_0_8 (.Z (\b[9] ), .A (B[9]), .B (n_0_8), .S (B[31]));
MUX2_X2 i_0_0_7 (.Z (\b[8] ), .A (B[8]), .B (n_0_7), .S (B[31]));
MUX2_X2 i_0_0_6 (.Z (\b[7] ), .A (B[7]), .B (n_0_6), .S (B[31]));
MUX2_X2 i_0_0_5 (.Z (\b[6] ), .A (B[6]), .B (n_0_5), .S (B[31]));
MUX2_X2 i_0_0_4 (.Z (spt__n6), .A (B[5]), .B (n_0_4), .S (B[31]));
MUX2_X2 i_0_0_3 (.Z (\b[4] ), .A (B[4]), .B (n_0_3), .S (B[31]));
MUX2_X2 i_0_0_2 (.Z (\b[3] ), .A (B[3]), .B (n_0_2), .S (B[31]));
MUX2_X2 i_0_0_1 (.Z (\b[2] ), .A (B[2]), .B (n_0_1), .S (B[31]));
MUX2_X1 i_0_0_0 (.Z (\b[1] ), .A (B[1]), .B (n_0_0), .S (B[31]));
WTM8__0_153 M14 (.Result ({\P[14][15] , \P[14][14] , \P[14][13] , \P[14][12] , \P[14][11] , 
    \P[14][10] , \P[14][9] , \P[14][8] , \P[14][7] , \P[14][6] , \P[14][5] , \P[14][4] , 
    \P[14][3] , \P[14][2] , \P[14][1] , \P[14][0] }), .A ({\a[31] , \a[30] , \a[29] , 
    \a[28] , \a[27] , \a[26] , \a[25] , \a[24] }), .B ({\b[23] , \b[22] , \b[21] , 
    \b[20] , \b[19] , \b[18] , \b[17] , \b[16] }));
adder64__0_154 A14 (.z ({\out[63] , \out[62] , \out[61] , \out[60] , \out[59] , \out[58] , 
    \out[57] , \out[56] , \out[55] , \out[54] , \out[53] , \out[52] , \out[51] , 
    \out[50] , \out[49] , \out[48] , \out[47] , \out[46] , \out[45] , \out[44] , 
    \out[43] , \out[42] , \out[41] , \out[40] , \out[39] , \out[38] , \out[37] , 
    \out[36] , \out[35] , \out[34] , \out[33] , \out[32] , \out[31] , \out[30] , 
    \out[29] , \out[28] , \out[27] , \out[26] , \out[25] , \out[24] , \out[23] , 
    \out[22] , \out[21] , \out[20] , \out[19] , \out[18] , \out[17] , \out[16] , 
    uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, uc_997, uc_998, 
    uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004}), .x ({uc_944, uc_945, uc_946, 
    uc_947, uc_948, uc_949, uc_950, uc_951, uc_952, uc_953, uc_954, uc_955, uc_956, 
    \Eight[0][50] , \Eight[0][49] , \Eight[0][48] , \Eight[0][47] , \Eight[0][46] , 
    \Eight[0][45] , \Eight[0][44] , \Eight[0][43] , \Eight[0][42] , \Eight[0][41] , 
    \Eight[0][40] , \Eight[0][39] , \Eight[0][38] , \Eight[0][37] , \Eight[0][36] , 
    \Eight[0][35] , \Eight[0][34] , \Eight[0][33] , \Eight[0][32] , \Eight[0][31] , 
    \Eight[0][30] , \Eight[0][29] , \Eight[0][28] , \Eight[0][27] , \Eight[0][26] , 
    \Eight[0][25] , \Eight[0][24] , \Eight[0][23] , \Eight[0][22] , \Eight[0][21] , 
    \Eight[0][20] , \Eight[0][19] , \Eight[0][18] , \Eight[0][17] , \Eight[0][16] , 
    uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, uc_963, uc_964, uc_965, uc_966, 
    uc_967, uc_968, uc_969, uc_970, uc_971, uc_972}), .y ({\Eight[1][63] , \Eight[1][62] , 
    \Eight[1][61] , \Eight[1][60] , \Eight[1][59] , \Eight[1][58] , \Eight[1][57] , 
    \Eight[1][56] , \Eight[1][55] , \Eight[1][54] , \Eight[1][53] , \Eight[1][52] , 
    \Eight[1][51] , \Eight[1][50] , \Eight[1][49] , \Eight[1][48] , \Eight[1][47] , 
    \Eight[1][46] , \Eight[1][45] , \Eight[1][44] , \Eight[1][43] , \Eight[1][42] , 
    \Eight[1][41] , \Eight[1][40] , \Eight[1][39] , \Eight[1][38] , \Eight[1][37] , 
    \Eight[1][36] , \Eight[1][35] , \Eight[1][34] , \Eight[1][33] , \Eight[1][32] , 
    \Eight[1][31] , \Eight[1][30] , \Eight[1][29] , \Eight[1][28] , \Eight[1][27] , 
    \Eight[1][26] , \Eight[1][25] , \Eight[1][24] , \Eight[1][23] , \Eight[1][22] , 
    \Eight[1][21] , \Eight[1][20] , \Eight[1][19] , \Eight[1][18] , \Eight[1][17] , 
    \Eight[1][16] , uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, uc_980, 
    uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, uc_987, uc_988}));
datapath i_0_6 (.p_0 ({n_0_62, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, 
    n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
    n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, 
    n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
    n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, 
    n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, 
    n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, uc_943}), .out ({
    \out[63] , \out[62] , \out[61] , \out[60] , \out[59] , \out[58] , \out[57] , 
    \out[56] , \out[55] , \out[54] , \out[53] , \out[52] , \out[51] , \out[50] , 
    \out[49] , \out[48] , \out[47] , \out[46] , \out[45] , \out[44] , \out[43] , 
    \out[42] , \out[41] , \out[40] , \out[39] , \out[38] , \out[37] , \out[36] , 
    \out[35] , \out[34] , \out[33] , \out[32] , \out[31] , \out[30] , \out[29] , 
    \out[28] , \out[27] , \out[26] , \out[25] , \out[24] , \out[23] , \out[22] , 
    \out[21] , \out[20] , \out[19] , \out[18] , \out[17] , \out[16] , \Eight[0][15] , 
    \Eight[0][14] , \Eight[0][13] , \Eight[0][12] , \Eight[0][11] , \Eight[0][10] , 
    \Eight[0][9] , \Eight[0][8] , \P[0][7] , \P[0][6] , \P[0][5] , \P[0][4] , \P[0][3] , 
    \P[0][2] , \P[0][1] , Result[0]}));
WTM8__1_2406 M10 (.Result ({\P[10][15] , \P[10][14] , \P[10][13] , \P[10][12] , \P[10][11] , 
    \P[10][10] , \P[10][9] , \P[10][8] , \P[10][7] , \P[10][6] , \P[10][5] , \P[10][4] , 
    \P[10][3] , \P[10][2] , \P[10][1] , \P[10][0] }), .A ({\a[23] , \a[22] , \a[21] , 
    \a[20] , \a[19] , \a[18] , \a[17] , \a[16] }), .B ({\b[23] , \b[22] , \b[21] , 
    \b[20] , \b[19] , \b[18] , \b[17] , \b[16] }), .A_5_PP_0 (spw__n50), .A_5_PP_1 (spw__n51)
    , .A_3_PP_0 (spw__n111), .A_4_PP_0 (spw__n122), .A_4_PP_1 (spw__n124));
datapath__0_79 i_0_3 (.p_0 ({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, 
    n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, 
    n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, 
    n_0_34, n_0_33, n_0_32, n_0_31, uc_942}), .A ({A[31], A[30], A[29], A[28], A[27], 
    A[26], A[25], A[24], A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], 
    A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
    A[3], A[2], A[1], A[0]}));
datapath__0_81 i_0_1 (.p_0 ({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
    n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
    n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
    n_0_2, n_0_1, n_0_0, uc_941}), .B ({B[31], B[30], B[29], B[28], B[27], B[26], 
    B[25], B[24], B[23], B[22], B[21], B[20], B[19], B[18], B[17], B[16], B[15], 
    B[14], B[13], B[12], B[11], B[10], B[9], B[8], B[7], B[6], B[5], B[4], B[3], 
    B[2], B[1], B[0]}));
adder64__1_3757 A12 (.z ({uc_920, uc_921, uc_922, uc_923, uc_924, uc_925, uc_926, 
    uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, \Eight[0][50] , \Eight[0][49] , 
    \Eight[0][48] , \Eight[0][47] , \Eight[0][46] , \Eight[0][45] , \Eight[0][44] , 
    \Eight[0][43] , \Eight[0][42] , \Eight[0][41] , \Eight[0][40] , \Eight[0][39] , 
    \Eight[0][38] , \Eight[0][37] , \Eight[0][36] , \Eight[0][35] , \Eight[0][34] , 
    \Eight[0][33] , \Eight[0][32] , \Eight[0][31] , \Eight[0][30] , \Eight[0][29] , 
    \Eight[0][28] , \Eight[0][27] , \Eight[0][26] , \Eight[0][25] , \Eight[0][24] , 
    \Eight[0][23] , \Eight[0][22] , \Eight[0][21] , \Eight[0][20] , \Eight[0][19] , 
    \Eight[0][18] , \Eight[0][17] , \Eight[0][16] , \Eight[0][15] , \Eight[0][14] , 
    \Eight[0][13] , \Eight[0][12] , \Eight[0][11] , \Eight[0][10] , \Eight[0][9] , 
    \Eight[0][8] , uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, uc_940})
    , .x ({uc_868, uc_869, uc_870, uc_871, uc_872, uc_873, uc_874, uc_875, uc_876, 
    uc_877, uc_878, uc_879, uc_880, uc_881, uc_882, uc_883, uc_884, uc_885, uc_886, 
    uc_887, uc_888, uc_889, \Quadruple[0][41] , \Quadruple[0][40] , \Quadruple[0][39] , 
    \Quadruple[0][38] , \Quadruple[0][37] , \Quadruple[0][36] , \Quadruple[0][35] , 
    \Quadruple[0][34] , \Quadruple[0][33] , \Quadruple[0][32] , \Quadruple[0][31] , 
    \Quadruple[0][30] , \Quadruple[0][29] , \Quadruple[0][28] , \Quadruple[0][27] , 
    \Quadruple[0][26] , \Quadruple[0][25] , \Quadruple[0][24] , \Quadruple[0][23] , 
    \Quadruple[0][22] , \Quadruple[0][21] , \Quadruple[0][20] , \Quadruple[0][19] , 
    \Quadruple[0][18] , \Quadruple[0][17] , \Quadruple[0][16] , \couple[0][15] , 
    \couple[0][14] , \couple[0][13] , \couple[0][12] , \couple[0][11] , \couple[0][10] , 
    \couple[0][9] , \couple[0][8] , uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, 
    uc_896, uc_897}), .y ({uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, 
    uc_905, uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, \Quadruple[1][49] , \Quadruple[1][48] , 
    \Quadruple[1][47] , \Quadruple[1][46] , \Quadruple[1][45] , \Quadruple[1][44] , 
    \Quadruple[1][43] , \Quadruple[1][42] , \Quadruple[1][41] , \Quadruple[1][40] , 
    \Quadruple[1][39] , \Quadruple[1][38] , \Quadruple[1][37] , \Quadruple[1][36] , 
    \Quadruple[1][35] , \Quadruple[1][34] , \Quadruple[1][33] , \Quadruple[1][32] , 
    \Quadruple[1][31] , \Quadruple[1][30] , \Quadruple[1][29] , \Quadruple[1][28] , 
    \Quadruple[1][27] , \Quadruple[1][26] , \Quadruple[1][25] , \Quadruple[1][24] , 
    \couple[2][23] , \couple[2][22] , \couple[2][21] , \couple[2][20] , \couple[2][19] , 
    \couple[2][18] , \couple[2][17] , \couple[2][16] , \P[4][7] , \P[4][6] , \P[4][5] , 
    \P[4][4] , \P[4][3] , \P[4][2] , \P[4][1] , \P[4][0] , uc_912, uc_913, uc_914, 
    uc_915, uc_916, uc_917, uc_918, uc_919}));
adder64__1_3564 A9 (.z ({uc_830, uc_831, uc_832, uc_833, uc_834, uc_835, uc_836, 
    uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, \Quadruple[1][49] , \Quadruple[1][48] , 
    \Quadruple[1][47] , \Quadruple[1][46] , \Quadruple[1][45] , \Quadruple[1][44] , 
    \Quadruple[1][43] , \Quadruple[1][42] , \Quadruple[1][41] , \Quadruple[1][40] , 
    \Quadruple[1][39] , \Quadruple[1][38] , \Quadruple[1][37] , \Quadruple[1][36] , 
    \Quadruple[1][35] , \Quadruple[1][34] , \Quadruple[1][33] , \Quadruple[1][32] , 
    \Quadruple[1][31] , \Quadruple[1][30] , \Quadruple[1][29] , \Quadruple[1][28] , 
    \Quadruple[1][27] , \Quadruple[1][26] , \Quadruple[1][25] , \Quadruple[1][24] , 
    uc_844, uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, uc_852, uc_853, 
    uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, uc_860, uc_861, uc_862, uc_863, 
    uc_864, uc_865, uc_866, uc_867}), .x ({uc_736, uc_737, uc_738, uc_739, uc_740, 
    uc_741, uc_742, uc_743, uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, 
    uc_751, uc_752, uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, uc_760, 
    uc_761, uc_762, uc_763, uc_764, uc_765, uc_766, \couple[2][32] , \couple[2][31] , 
    \couple[2][30] , \couple[2][29] , \couple[2][28] , \couple[2][27] , \couple[2][26] , 
    \couple[2][25] , \couple[2][24] , uc_767, uc_768, uc_769, uc_770, uc_771, uc_772, 
    uc_773, uc_774, uc_775, uc_776, uc_777, uc_778, uc_779, uc_780, uc_781, uc_782, 
    uc_783, uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, uc_790}), .y ({uc_791, 
    uc_792, uc_793, uc_794, uc_795, uc_796, uc_797, uc_798, uc_799, uc_800, uc_801, 
    uc_802, uc_803, uc_804, uc_805, \couple[3][48] , \couple[3][47] , \couple[3][46] , 
    \couple[3][45] , \couple[3][44] , \couple[3][43] , \couple[3][42] , \couple[3][41] , 
    \couple[3][40] , \couple[3][39] , \couple[3][38] , \couple[3][37] , \couple[3][36] , 
    \couple[3][35] , \couple[3][34] , \couple[3][33] , \couple[3][32] , \P[6][7] , 
    \P[6][6] , \P[6][5] , \P[6][4] , \P[6][3] , \P[6][2] , \P[6][1] , \P[6][0] , 
    uc_806, uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, 
    uc_816, uc_817, uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, 
    uc_826, uc_827, uc_828, uc_829}));
adder64__1_3371 A3 (.z ({uc_689, uc_690, uc_691, uc_692, uc_693, uc_694, uc_695, 
    uc_696, uc_697, uc_698, uc_699, uc_700, uc_701, uc_702, uc_703, \couple[3][48] , 
    \couple[3][47] , \couple[3][46] , \couple[3][45] , \couple[3][44] , \couple[3][43] , 
    \couple[3][42] , \couple[3][41] , \couple[3][40] , \couple[3][39] , \couple[3][38] , 
    \couple[3][37] , \couple[3][36] , \couple[3][35] , \couple[3][34] , \couple[3][33] , 
    \couple[3][32] , uc_704, uc_705, uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, 
    uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, uc_719, uc_720, uc_721, 
    uc_722, uc_723, uc_724, uc_725, uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, 
    uc_732, uc_733, uc_734, uc_735}), .x ({uc_585, uc_586, uc_587, uc_588, uc_589, 
    uc_590, uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, 
    uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, uc_607, uc_608, \P[6][15] , 
    \P[6][14] , \P[6][13] , \P[6][12] , \P[6][11] , \P[6][10] , \P[6][9] , \P[6][8] , 
    uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, uc_616, uc_617, uc_618, 
    uc_619, uc_620, uc_621, uc_622, uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, 
    uc_629, uc_630, uc_631, uc_632, uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, 
    uc_639, uc_640}), .y ({uc_641, uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, 
    uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, uc_654, uc_655, uc_656, \P[7][15] , 
    \P[7][14] , \P[7][13] , \P[7][12] , \P[7][11] , \P[7][10] , \P[7][9] , \P[7][8] , 
    \P[7][7] , \P[7][6] , \P[7][5] , \P[7][4] , \P[7][3] , \P[7][2] , \P[7][1] , 
    \P[7][0] , uc_657, uc_658, uc_659, uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, 
    uc_666, uc_667, uc_668, uc_669, uc_670, uc_671, uc_672, uc_673, uc_674, uc_675, 
    uc_676, uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, 
    uc_686, uc_687, uc_688}));
WTM8__1_2152 M7 (.Result ({\P[7][15] , \P[7][14] , \P[7][13] , \P[7][12] , \P[7][11] , 
    \P[7][10] , \P[7][9] , \P[7][8] , \P[7][7] , \P[7][6] , \P[7][5] , \P[7][4] , 
    \P[7][3] , \P[7][2] , \P[7][1] , \P[7][0] }), .A ({\a[15] , \a[14] , \a[13] , 
    \a[12] , \a[11] , \a[10] , \a[9] , \a[8] }), .B ({\b[31] , \b[30] , \b[29] , 
    \b[28] , \b[27] , \b[26] , \b[25] , \b[24] }), .A_7_PP_0 (\a[15] ));
WTM8__1_1898 M6 (.Result ({\P[6][15] , \P[6][14] , \P[6][13] , \P[6][12] , \P[6][11] , 
    \P[6][10] , \P[6][9] , \P[6][8] , \P[6][7] , \P[6][6] , \P[6][5] , \P[6][4] , 
    \P[6][3] , \P[6][2] , \P[6][1] , \P[6][0] }), .A ({\a[15] , \a[14] , \a[13] , 
    \a[12] , \a[11] , \a[10] , \a[9] , \a[8] }), .B ({\b[23] , \b[22] , \b[21] , 
    \b[20] , \b[19] , \b[18] , \b[17] , \b[16] }), .A_5_PP_0 (spw__n80), .A_6_PP_0 (spw__n166)
    , .A_7_PP_0 (spw__n182), .A_7_PP_1 (spw__n183));
adder64__1_3178 A2 (.z ({uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, 
    uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, 
    uc_555, uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, 
    uc_565, uc_566, uc_567, uc_568, \couple[2][32] , \couple[2][31] , \couple[2][30] , 
    \couple[2][29] , \couple[2][28] , \couple[2][27] , \couple[2][26] , \couple[2][25] , 
    \couple[2][24] , \couple[2][23] , \couple[2][22] , \couple[2][21] , \couple[2][20] , 
    \couple[2][19] , \couple[2][18] , \couple[2][17] , \couple[2][16] , uc_569, uc_570, 
    uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, uc_580, 
    uc_581, uc_582, uc_583, uc_584}), .x ({uc_434, uc_435, uc_436, uc_437, uc_438, 
    uc_439, uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, 
    uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, 
    uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, 
    uc_469, uc_470, uc_471, uc_472, uc_473, \P[4][15] , \P[4][14] , \P[4][13] , \P[4][12] , 
    \P[4][11] , \P[4][10] , \P[4][9] , \P[4][8] , uc_474, uc_475, uc_476, uc_477, 
    uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, 
    uc_488, uc_489}), .y ({uc_490, uc_491, uc_492, uc_493, uc_494, uc_495, uc_496, 
    uc_497, uc_498, uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, 
    uc_507, uc_508, uc_509, uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, 
    uc_517, uc_518, uc_519, uc_520, uc_521, \P[5][15] , \P[5][14] , \P[5][13] , \P[5][12] , 
    \P[5][11] , \P[5][10] , \P[5][9] , \P[5][8] , \P[5][7] , \P[5][6] , \P[5][5] , 
    \P[5][4] , \P[5][3] , \P[5][2] , \P[5][1] , \P[5][0] , uc_522, uc_523, uc_524, 
    uc_525, uc_526, uc_527, uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, 
    uc_535, uc_536, uc_537}));
WTM8__1_1644 M5 (.Result ({\P[5][15] , \P[5][14] , \P[5][13] , \P[5][12] , \P[5][11] , 
    \P[5][10] , \P[5][9] , \P[5][8] , \P[5][7] , \P[5][6] , \P[5][5] , \P[5][4] , 
    \P[5][3] , \P[5][2] , \P[5][1] , \P[5][0] }), .A ({spw__n183, spw__n166, spw__n80, 
    \a[12] , \a[11] , \a[10] , \a[9] , \a[8] }), .B ({\b[15] , \b[14] , spw__n226, 
    \b[12] , \b[11] , \b[10] , \b[9] , \b[8] }), .B_7_PP_0 (\b[15] ), .B_5_PP_0 (spw__n226));
WTM8__1_1390 M4 (.Result ({\P[4][15] , \P[4][14] , \P[4][13] , \P[4][12] , \P[4][11] , 
    \P[4][10] , \P[4][9] , \P[4][8] , \P[4][7] , \P[4][6] , \P[4][5] , \P[4][4] , 
    \P[4][3] , \P[4][2] , \P[4][1] , \P[4][0] }), .A ({spw__n183, spw__n166, spw__n80, 
    \a[12] , \a[11] , \a[10] , \a[9] , \a[8] }), .B ({\b[7] , \b[6] , \b[5] , \b[4] , 
    \b[3] , \b[2] , \b[1] , B[0]}));
adder64__1_2985 A8 (.z ({uc_396, uc_397, uc_398, uc_399, uc_400, uc_401, uc_402, 
    uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, uc_409, uc_410, uc_411, uc_412, 
    uc_413, uc_414, uc_415, uc_416, uc_417, \Quadruple[0][41] , \Quadruple[0][40] , 
    \Quadruple[0][39] , \Quadruple[0][38] , \Quadruple[0][37] , \Quadruple[0][36] , 
    \Quadruple[0][35] , \Quadruple[0][34] , \Quadruple[0][33] , \Quadruple[0][32] , 
    \Quadruple[0][31] , \Quadruple[0][30] , \Quadruple[0][29] , \Quadruple[0][28] , 
    \Quadruple[0][27] , \Quadruple[0][26] , \Quadruple[0][25] , \Quadruple[0][24] , 
    \Quadruple[0][23] , \Quadruple[0][22] , \Quadruple[0][21] , \Quadruple[0][20] , 
    \Quadruple[0][19] , \Quadruple[0][18] , \Quadruple[0][17] , \Quadruple[0][16] , 
    uc_418, uc_419, uc_420, uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, 
    uc_428, uc_429, uc_430, uc_431, uc_432, uc_433}), .x ({uc_302, uc_303, uc_304, 
    uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, uc_313, uc_314, 
    uc_315, uc_316, uc_317, uc_318, uc_319, uc_320, uc_321, uc_322, uc_323, uc_324, 
    uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, uc_334, 
    uc_335, uc_336, uc_337, uc_338, uc_339, uc_340, \couple[0][24] , \couple[0][23] , 
    \couple[0][22] , \couple[0][21] , \couple[0][20] , \couple[0][19] , \couple[0][18] , 
    \couple[0][17] , \couple[0][16] , uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, 
    uc_347, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356})
    , .y ({uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, 
    uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, 
    uc_376, uc_377, uc_378, uc_379, \couple[1][40] , \couple[1][39] , \couple[1][38] , 
    \couple[1][37] , \couple[1][36] , \couple[1][35] , \couple[1][34] , \couple[1][33] , 
    \couple[1][32] , \couple[1][31] , \couple[1][30] , \couple[1][29] , \couple[1][28] , 
    \couple[1][27] , \couple[1][26] , \couple[1][25] , \couple[1][24] , \P[2][7] , 
    \P[2][6] , \P[2][5] , \P[2][4] , \P[2][3] , \P[2][2] , \P[2][1] , \P[2][0] , 
    uc_380, uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, 
    uc_390, uc_391, uc_392, uc_393, uc_394, uc_395}));
adder64__1_2792 A1 (.z ({uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, 
    uc_262, uc_263, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, 
    uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, \couple[1][40] , \couple[1][39] , 
    \couple[1][38] , \couple[1][37] , \couple[1][36] , \couple[1][35] , \couple[1][34] , 
    \couple[1][33] , \couple[1][32] , \couple[1][31] , \couple[1][30] , \couple[1][29] , 
    \couple[1][28] , \couple[1][27] , \couple[1][26] , \couple[1][25] , \couple[1][24] , 
    uc_278, uc_279, uc_280, uc_281, uc_282, uc_283, uc_284, uc_285, uc_286, uc_287, 
    uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297, 
    uc_298, uc_299, uc_300, uc_301}), .x ({uc_151, uc_152, uc_153, uc_154, uc_155, 
    uc_156, uc_157, uc_158, uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, 
    uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, 
    uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, \P[2][15] , \P[2][14] , 
    \P[2][13] , \P[2][12] , \P[2][11] , \P[2][10] , \P[2][9] , \P[2][8] , uc_183, 
    uc_184, uc_185, uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192, uc_193, 
    uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, 
    uc_204, uc_205, uc_206}), .y ({uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, 
    uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, 
    uc_223, uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, \P[3][15] , \P[3][14] , 
    \P[3][13] , \P[3][12] , \P[3][11] , \P[3][10] , \P[3][9] , \P[3][8] , \P[3][7] , 
    \P[3][6] , \P[3][5] , \P[3][4] , \P[3][3] , \P[3][2] , \P[3][1] , \P[3][0] , 
    uc_231, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, uc_239, uc_240, 
    uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, uc_248, uc_249, uc_250, 
    uc_251, uc_252, uc_253, uc_254}));
WTM8__1_1136 M3 (.Result ({\P[3][15] , \P[3][14] , \P[3][13] , \P[3][12] , \P[3][11] , 
    \P[3][10] , \P[3][9] , \P[3][8] , \P[3][7] , \P[3][6] , \P[3][5] , \P[3][4] , 
    \P[3][3] , \P[3][2] , \P[3][1] , \P[3][0] }), .A ({\a[7] , \a[6] , \a[5] , \a[4] , 
    \a[3] , \a[2] , \a[1] , A[0]}), .B ({\b[31] , \b[30] , \b[29] , \b[28] , \b[27] , 
    \b[26] , \b[25] , \b[24] }));
WTM8__1_882 M2 (.Result ({\P[2][15] , \P[2][14] , \P[2][13] , \P[2][12] , \P[2][11] , 
    \P[2][10] , \P[2][9] , \P[2][8] , \P[2][7] , \P[2][6] , \P[2][5] , \P[2][4] , 
    \P[2][3] , \P[2][2] , \P[2][1] , \P[2][0] }), .A ({\a[7] , \a[6] , \a[5] , \a[4] , 
    \a[3] , \a[2] , \a[1] , A[0]}), .B ({\b[23] , \b[22] , \b[21] , \b[20] , \b[19] , 
    \b[18] , \b[17] , \b[16] }), .A_7_PP_0 (spw__n67), .A_6_PP_0 (spw__n276), .A_5_PP_0 (spw__n88)
    , .A_5_PP_1 (spw__n89), .A_6_PP_0PP_0 (spw__n277));
adder64__1_2599 A0 (.z ({uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, 
    uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, 
    uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, uc_127, uc_128, uc_129, uc_130, 
    uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, 
    uc_141, uc_142, \couple[0][24] , \couple[0][23] , \couple[0][22] , \couple[0][21] , 
    \couple[0][20] , \couple[0][19] , \couple[0][18] , \couple[0][17] , \couple[0][16] , 
    \couple[0][15] , \couple[0][14] , \couple[0][13] , \couple[0][12] , \couple[0][11] , 
    \couple[0][10] , \couple[0][9] , \couple[0][8] , uc_143, uc_144, uc_145, uc_146, 
    uc_147, uc_148, uc_149, uc_150}), .x ({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
    uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, 
    uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, 
    uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, 
    uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, \P[0][15] , \P[0][14] , \P[0][13] , 
    \P[0][12] , \P[0][11] , \P[0][10] , \P[0][9] , \P[0][8] , uc_48, uc_49, uc_50, 
    uc_51, uc_52, uc_53, uc_54, uc_55}), .y ({uc_56, uc_57, uc_58, uc_59, uc_60, 
    uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, 
    uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, 
    uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
    uc_94, uc_95, \P[1][15] , \P[1][14] , \P[1][13] , \P[1][12] , \P[1][11] , \P[1][10] , 
    \P[1][9] , \P[1][8] , \P[1][7] , \P[1][6] , \P[1][5] , \P[1][4] , \P[1][3] , 
    \P[1][2] , \P[1][1] , \P[1][0] , uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, 
    uc_102, uc_103}));
WTM8__1_628 M0 (.Result ({\P[0][15] , \P[0][14] , \P[0][13] , \P[0][12] , \P[0][11] , 
    \P[0][10] , \P[0][9] , \P[0][8] , \P[0][7] , \P[0][6] , \P[0][5] , \P[0][4] , 
    \P[0][3] , \P[0][2] , \P[0][1] , Result[0]}), .A ({spw__n325, spw__n277, spw__n90, 
    \a[4] , \a[3] , \a[2] , \a[1] , A[0]}), .B ({\b[7] , \b[6] , \b[5] , \b[4] , 
    \b[3] , \b[2] , \b[1] , B[0]}), .B_5_PP_0 (spw__n314));
CLKBUF_X3 sps__L1_c1 (.Z (sps__n1), .A (n_0_0_0));
BUF_X4 spt__c6 (.Z (spw__n314), .A (spt__n6));
BUF_X4 spw__c259 (.Z (\a[18] ), .A (spw__n384));
BUF_X4 spt__c12 (.Z (spw__n90), .A (spt__n12));
BUF_X1 spw__L3_c3_c34 (.Z (\a[21] ), .A (spw__n50));
BUF_X2 spw__L2_c2_c35 (.Z (spw__n50), .A (spw__n51));
BUF_X1 spw__L1_c1_c36 (.Z (spw__n51), .A (spw__n54));
BUF_X4 spw__L2_c6_c37 (.Z (spw__n52), .A (spw__n53));
BUF_X1 spw__L1_c5_c38 (.Z (spw__n53), .A (spw__n54));
BUF_X4 spw__L2_c2_c51 (.Z (\a[7] ), .A (spw__n67));
BUF_X4 spw__L1_c1_c52 (.Z (spw__n67), .A (spt__n3));
BUF_X4 spw__L1_c1_c59 (.Z (\a[6] ), .A (spt__n9));
BUF_X2 spw__L2_c2_c64 (.Z (\a[13] ), .A (spw__n80));
BUF_X4 spw__L1_c1_c65 (.Z (spw__n80), .A (spw__n81));
BUF_X4 spw__L3_c3_c72 (.Z (\a[5] ), .A (spw__n88));
BUF_X2 spw__L2_c2_c73 (.Z (spw__n88), .A (spw__n89));
BUF_X1 spw__L1_c1_c74 (.Z (spw__n89), .A (spw__n90));
BUF_X1 spw__L3_c3_c85 (.Z (\a[19] ), .A (spw__n111));
BUF_X2 spw__L2_c2_c86 (.Z (spw__n111), .A (spw__n112));
BUF_X4 spw__L1_c1_c87 (.Z (spw__n112), .A (spw__n113));
BUF_X4 spw__L2_c2_c96 (.Z (\a[20] ), .A (spw__n122));
BUF_X1 spw__L1_c1_c97 (.Z (spw__n122), .A (spw__n124));
BUF_X1 spw__L1_c4_c98 (.Z (spw__n123), .A (spw__n124));
BUF_X2 spw__L3_c3_c107 (.Z (\b[15] ), .A (spw__n135));
BUF_X2 spw__L2_c2_c108 (.Z (spw__n135), .A (spw__n136));
BUF_X1 spw__L1_c1_c109 (.Z (spw__n136), .A (spw__n139));
BUF_X1 spw__L2_c6_c110 (.Z (spw__n137), .A (spw__n138));
BUF_X2 spw__L1_c5_c111 (.Z (spw__n138), .A (spw__n139));
BUF_X4 spw__L4_c4_c124 (.Z (\a[22] ), .A (spw__n152));
BUF_X1 spw__L3_c3_c125 (.Z (spw__n152), .A (spw__n153));
BUF_X2 spw__L2_c2_c126 (.Z (spw__n153), .A (spw__n154));
BUF_X1 spw__L1_c1_c127 (.Z (spw__n154), .A (spw__n155));
BUF_X4 spw__L2_c2_c138 (.Z (\a[14] ), .A (spw__n166));
BUF_X4 spw__L1_c1_c139 (.Z (spw__n166), .A (spw__n167));
BUF_X2 spw__L3_c3_c146 (.Z (\a[15] ), .A (spw__n182));
BUF_X1 spw__L2_c2_c147 (.Z (spw__n182), .A (spw__n183));
BUF_X4 spw__L1_c1_c148 (.Z (spw__n183), .A (spw__n184));
BUF_X4 spw__L2_c2_c161 (.Z (\a[23] ), .A (spw__n215));
BUF_X1 spw__L1_c1_c162 (.Z (spw__n215), .A (spw__n216));
BUF_X2 spw__L2_c2_c169 (.Z (\b[13] ), .A (spw__n225));
BUF_X2 spw__L1_c1_c170 (.Z (spw__n225), .A (spw__n230));
BUF_X2 spw__L4_c7_c171 (.Z (spw__n226), .A (spw__n227));
BUF_X1 spw__L3_c6_c172 (.Z (spw__n227), .A (spw__n228));
BUF_X1 spw__L2_c5_c173 (.Z (spw__n228), .A (spw__n229));
BUF_X2 spw__L1_c4_c174 (.Z (spw__n229), .A (spw__n230));
BUF_X4 spw__L1_c1_c223 (.Z (\b[5] ), .A (spw__n314));
BUF_X1 spw__L3_c3_c206 (.Z (spt__n9), .A (spw__n276));
BUF_X1 spw__L2_c2_c207 (.Z (spw__n276), .A (spw__n277));
BUF_X8 spw__L1_c1_c208 (.Z (spw__n277), .A (spw__n278));
CLKBUF_X1 spw__L2_c2_c233 (.Z (spt__n3), .A (spw__n324));
CLKBUF_X1 spw__L1_c1_c234 (.Z (spw__n324), .A (spw__n325));

endmodule //WTM32

module registered_WTM (A, B, Result, clk, reset);

output [63:0] Result;
input [31:0] A;
input [31:0] B;
input clk;
input reset;
wire \Result_OUT[63] ;
wire \Result_OUT[62] ;
wire \Result_OUT[61] ;
wire \Result_OUT[60] ;
wire \Result_OUT[59] ;
wire \Result_OUT[58] ;
wire \Result_OUT[57] ;
wire \Result_OUT[56] ;
wire \Result_OUT[55] ;
wire \Result_OUT[54] ;
wire \Result_OUT[53] ;
wire \Result_OUT[52] ;
wire \Result_OUT[51] ;
wire \Result_OUT[50] ;
wire \Result_OUT[49] ;
wire \Result_OUT[48] ;
wire \Result_OUT[47] ;
wire \Result_OUT[46] ;
wire \Result_OUT[45] ;
wire \Result_OUT[44] ;
wire \Result_OUT[43] ;
wire \Result_OUT[42] ;
wire \Result_OUT[41] ;
wire \Result_OUT[40] ;
wire \Result_OUT[39] ;
wire \Result_OUT[38] ;
wire \Result_OUT[37] ;
wire \Result_OUT[36] ;
wire \Result_OUT[35] ;
wire \Result_OUT[34] ;
wire \Result_OUT[33] ;
wire \Result_OUT[32] ;
wire \Result_OUT[31] ;
wire \Result_OUT[30] ;
wire \Result_OUT[29] ;
wire \Result_OUT[28] ;
wire \Result_OUT[27] ;
wire \Result_OUT[26] ;
wire \Result_OUT[25] ;
wire \Result_OUT[24] ;
wire \Result_OUT[23] ;
wire \Result_OUT[22] ;
wire \Result_OUT[21] ;
wire \Result_OUT[20] ;
wire \Result_OUT[19] ;
wire \Result_OUT[18] ;
wire \Result_OUT[17] ;
wire \Result_OUT[16] ;
wire \Result_OUT[15] ;
wire \Result_OUT[14] ;
wire \Result_OUT[13] ;
wire \Result_OUT[12] ;
wire \Result_OUT[11] ;
wire \Result_OUT[10] ;
wire \Result_OUT[9] ;
wire \Result_OUT[8] ;
wire \Result_OUT[7] ;
wire \Result_OUT[6] ;
wire \Result_OUT[5] ;
wire \Result_OUT[4] ;
wire \Result_OUT[3] ;
wire \Result_OUT[2] ;
wire \Result_OUT[1] ;
wire \Result_OUT[0] ;
wire \A_IN[31] ;
wire \A_IN[30] ;
wire \A_IN[29] ;
wire \A_IN[28] ;
wire \A_IN[27] ;
wire \A_IN[26] ;
wire \A_IN[25] ;
wire \A_IN[24] ;
wire \A_IN[23] ;
wire \A_IN[22] ;
wire \A_IN[21] ;
wire \A_IN[20] ;
wire \A_IN[19] ;
wire \A_IN[18] ;
wire \A_IN[17] ;
wire \A_IN[16] ;
wire \A_IN[15] ;
wire \A_IN[14] ;
wire \A_IN[13] ;
wire \A_IN[12] ;
wire \A_IN[11] ;
wire \A_IN[10] ;
wire \A_IN[9] ;
wire \A_IN[8] ;
wire \A_IN[7] ;
wire \A_IN[6] ;
wire \A_IN[5] ;
wire \A_IN[4] ;
wire \A_IN[3] ;
wire \A_IN[2] ;
wire \A_IN[1] ;
wire \A_IN[0] ;
wire \B_IN[31] ;
wire \B_IN[30] ;
wire \B_IN[29] ;
wire \B_IN[28] ;
wire \B_IN[27] ;
wire \B_IN[26] ;
wire \B_IN[25] ;
wire \B_IN[24] ;
wire \B_IN[23] ;
wire \B_IN[22] ;
wire \B_IN[21] ;
wire \B_IN[20] ;
wire \B_IN[19] ;
wire \B_IN[18] ;
wire \B_IN[17] ;
wire \B_IN[16] ;
wire \B_IN[15] ;
wire \B_IN[14] ;
wire \B_IN[13] ;
wire \B_IN[12] ;
wire \B_IN[11] ;
wire \B_IN[10] ;
wire \B_IN[9] ;
wire \B_IN[8] ;
wire \B_IN[7] ;
wire \B_IN[6] ;
wire \B_IN[5] ;
wire \B_IN[4] ;
wire \B_IN[3] ;
wire \B_IN[2] ;
wire \B_IN[1] ;
wire \B_IN[0] ;


register__parameterized0 outputReg (.DATA_OUT ({Result[63], Result[62], Result[61], 
    Result[60], Result[59], Result[58], Result[57], Result[56], Result[55], Result[54], 
    Result[53], Result[52], Result[51], Result[50], Result[49], Result[48], Result[47], 
    Result[46], Result[45], Result[44], Result[43], Result[42], Result[41], Result[40], 
    Result[39], Result[38], Result[37], Result[36], Result[35], Result[34], Result[33], 
    Result[32], Result[31], Result[30], Result[29], Result[28], Result[27], Result[26], 
    Result[25], Result[24], Result[23], Result[22], Result[21], Result[20], Result[19], 
    Result[18], Result[17], Result[16], Result[15], Result[14], Result[13], Result[12], 
    Result[11], Result[10], Result[9], Result[8], Result[7], Result[6], Result[5], 
    Result[4], Result[3], Result[2], Result[1], Result[0]}), .DATA_IN ({\Result_OUT[63] , 
    \Result_OUT[62] , \Result_OUT[61] , \Result_OUT[60] , \Result_OUT[59] , \Result_OUT[58] , 
    \Result_OUT[57] , \Result_OUT[56] , \Result_OUT[55] , \Result_OUT[54] , \Result_OUT[53] , 
    \Result_OUT[52] , \Result_OUT[51] , \Result_OUT[50] , \Result_OUT[49] , \Result_OUT[48] , 
    \Result_OUT[47] , \Result_OUT[46] , \Result_OUT[45] , \Result_OUT[44] , \Result_OUT[43] , 
    \Result_OUT[42] , \Result_OUT[41] , \Result_OUT[40] , \Result_OUT[39] , \Result_OUT[38] , 
    \Result_OUT[37] , \Result_OUT[36] , \Result_OUT[35] , \Result_OUT[34] , \Result_OUT[33] , 
    \Result_OUT[32] , \Result_OUT[31] , \Result_OUT[30] , \Result_OUT[29] , \Result_OUT[28] , 
    \Result_OUT[27] , \Result_OUT[26] , \Result_OUT[25] , \Result_OUT[24] , \Result_OUT[23] , 
    \Result_OUT[22] , \Result_OUT[21] , \Result_OUT[20] , \Result_OUT[19] , \Result_OUT[18] , 
    \Result_OUT[17] , \Result_OUT[16] , \Result_OUT[15] , \Result_OUT[14] , \Result_OUT[13] , 
    \Result_OUT[12] , \Result_OUT[11] , \Result_OUT[10] , \Result_OUT[9] , \Result_OUT[8] , 
    \Result_OUT[7] , \Result_OUT[6] , \Result_OUT[5] , \Result_OUT[4] , \Result_OUT[3] , 
    \Result_OUT[2] , \Result_OUT[1] , \Result_OUT[0] }), .clk (clk), .reset (reset));
register inputReg_2 (.DATA_OUT ({\B_IN[31] , \B_IN[30] , \B_IN[29] , \B_IN[28] , 
    \B_IN[27] , \B_IN[26] , \B_IN[25] , \B_IN[24] , \B_IN[23] , \B_IN[22] , \B_IN[21] , 
    \B_IN[20] , \B_IN[19] , \B_IN[18] , \B_IN[17] , \B_IN[16] , \B_IN[15] , \B_IN[14] , 
    \B_IN[13] , \B_IN[12] , \B_IN[11] , \B_IN[10] , \B_IN[9] , \B_IN[8] , \B_IN[7] , 
    \B_IN[6] , \B_IN[5] , \B_IN[4] , \B_IN[3] , \B_IN[2] , \B_IN[1] , \B_IN[0] })
    , .DATA_IN ({B[31], B[30], B[29], B[28], B[27], B[26], B[25], B[24], B[23], B[22], 
    B[21], B[20], B[19], B[18], B[17], B[16], B[15], B[14], B[13], B[12], B[11], 
    B[10], B[9], B[8], B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .clk (clk), .reset (reset));
register__3_1 inputReg_1 (.DATA_OUT ({\A_IN[31] , \A_IN[30] , \A_IN[29] , \A_IN[28] , 
    \A_IN[27] , \A_IN[26] , \A_IN[25] , \A_IN[24] , \A_IN[23] , \A_IN[22] , \A_IN[21] , 
    \A_IN[20] , \A_IN[19] , \A_IN[18] , \A_IN[17] , \A_IN[16] , \A_IN[15] , \A_IN[14] , 
    \A_IN[13] , \A_IN[12] , \A_IN[11] , \A_IN[10] , \A_IN[9] , \A_IN[8] , \A_IN[7] , 
    \A_IN[6] , \A_IN[5] , \A_IN[4] , \A_IN[3] , \A_IN[2] , \A_IN[1] , \A_IN[0] })
    , .DATA_IN ({A[31], A[30], A[29], A[28], A[27], A[26], A[25], A[24], A[23], A[22], 
    A[21], A[20], A[19], A[18], A[17], A[16], A[15], A[14], A[13], A[12], A[11], 
    A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0]}), .clk (clk), .reset (reset));
WTM32 multiplier (.Result ({\Result_OUT[63] , \Result_OUT[62] , \Result_OUT[61] , 
    \Result_OUT[60] , \Result_OUT[59] , \Result_OUT[58] , \Result_OUT[57] , \Result_OUT[56] , 
    \Result_OUT[55] , \Result_OUT[54] , \Result_OUT[53] , \Result_OUT[52] , \Result_OUT[51] , 
    \Result_OUT[50] , \Result_OUT[49] , \Result_OUT[48] , \Result_OUT[47] , \Result_OUT[46] , 
    \Result_OUT[45] , \Result_OUT[44] , \Result_OUT[43] , \Result_OUT[42] , \Result_OUT[41] , 
    \Result_OUT[40] , \Result_OUT[39] , \Result_OUT[38] , \Result_OUT[37] , \Result_OUT[36] , 
    \Result_OUT[35] , \Result_OUT[34] , \Result_OUT[33] , \Result_OUT[32] , \Result_OUT[31] , 
    \Result_OUT[30] , \Result_OUT[29] , \Result_OUT[28] , \Result_OUT[27] , \Result_OUT[26] , 
    \Result_OUT[25] , \Result_OUT[24] , \Result_OUT[23] , \Result_OUT[22] , \Result_OUT[21] , 
    \Result_OUT[20] , \Result_OUT[19] , \Result_OUT[18] , \Result_OUT[17] , \Result_OUT[16] , 
    \Result_OUT[15] , \Result_OUT[14] , \Result_OUT[13] , \Result_OUT[12] , \Result_OUT[11] , 
    \Result_OUT[10] , \Result_OUT[9] , \Result_OUT[8] , \Result_OUT[7] , \Result_OUT[6] , 
    \Result_OUT[5] , \Result_OUT[4] , \Result_OUT[3] , \Result_OUT[2] , \Result_OUT[1] , 
    \Result_OUT[0] }), .A ({\A_IN[31] , \A_IN[30] , \A_IN[29] , \A_IN[28] , \A_IN[27] , 
    \A_IN[26] , \A_IN[25] , \A_IN[24] , \A_IN[23] , \A_IN[22] , \A_IN[21] , \A_IN[20] , 
    \A_IN[19] , \A_IN[18] , \A_IN[17] , \A_IN[16] , \A_IN[15] , \A_IN[14] , \A_IN[13] , 
    \A_IN[12] , \A_IN[11] , \A_IN[10] , \A_IN[9] , \A_IN[8] , \A_IN[7] , \A_IN[6] , 
    \A_IN[5] , \A_IN[4] , \A_IN[3] , \A_IN[2] , \A_IN[1] , \A_IN[0] }), .B ({\B_IN[31] , 
    \B_IN[30] , \B_IN[29] , \B_IN[28] , \B_IN[27] , \B_IN[26] , \B_IN[25] , \B_IN[24] , 
    \B_IN[23] , \B_IN[22] , \B_IN[21] , \B_IN[20] , \B_IN[19] , \B_IN[18] , \B_IN[17] , 
    \B_IN[16] , \B_IN[15] , \B_IN[14] , \B_IN[13] , \B_IN[12] , \B_IN[11] , \B_IN[10] , 
    \B_IN[9] , \B_IN[8] , \B_IN[7] , \B_IN[6] , \B_IN[5] , \B_IN[4] , \B_IN[3] , 
    \B_IN[2] , \B_IN[1] , \B_IN[0] }));

endmodule //registered_WTM


