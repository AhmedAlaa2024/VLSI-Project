/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Dec 24 01:25:08 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2636546320 */

module FA__1_627(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_624(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_621(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_615(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_612(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_609(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_606(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_603(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_600(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_597(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_594(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_591(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_588(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_585(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_582(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_579(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_576(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_573(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_567(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_564(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_561(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_558(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_555(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_552(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_549(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_546(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_543(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_540(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_537(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_534(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_531(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_528(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_525(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_519(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_516(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_513(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_510(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_507(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_504(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_501(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_495(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_492(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_489(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_486(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_483(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_480(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_477(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_474(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_471(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_468(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_465(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_462(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_459(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_456(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_453(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_447(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_444(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_441(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_628(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_627 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_624 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_621 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_618 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_615 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_612 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_609 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_606 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_603 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_600 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_597 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_594 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_591 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_588 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_585 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_582 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_579 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_576 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_573 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_570 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_567 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_564 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_561 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_558 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_555 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_552 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_549 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_546 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_543 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_540 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_537 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_534 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_531 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_528 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_525 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_522 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_519 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_516 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_513 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_510 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_507 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_504 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_501 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_498 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_495 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_492 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_489 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_486 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_483 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_480 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_477 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_474 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_471 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_468 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_465 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_462 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_459 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_456 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_453 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_450 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_447 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_444 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_441 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_2574(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_2571(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2568(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2565(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2559(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2556(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2553(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2550(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2547(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2544(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2541(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2538(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2535(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2532(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2529(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_2599(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_2574 genblk1_8_F (.a(x[8]), .b(y[8]), .cin(), .sum(z[8]), .carry(
      carry[8]));
   FA__1_2571 genblk1_9_F (.a(x[9]), .b(y[9]), .cin(carry[8]), .sum(z[9]), 
      .carry(carry[9]));
   FA__1_2568 genblk1_10_F (.a(x[10]), .b(y[10]), .cin(carry[9]), .sum(z[10]), 
      .carry(carry[10]));
   FA__1_2565 genblk1_11_F (.a(x[11]), .b(y[11]), .cin(carry[10]), .sum(z[11]), 
      .carry(carry[11]));
   FA__1_2562 genblk1_12_F (.a(x[12]), .b(y[12]), .cin(carry[11]), .sum(z[12]), 
      .carry(carry[12]));
   FA__1_2559 genblk1_13_F (.a(x[13]), .b(y[13]), .cin(carry[12]), .sum(z[13]), 
      .carry(carry[13]));
   FA__1_2556 genblk1_14_F (.a(x[14]), .b(y[14]), .cin(carry[13]), .sum(z[14]), 
      .carry(carry[14]));
   FA__1_2553 genblk1_15_F (.a(x[15]), .b(y[15]), .cin(carry[14]), .sum(z[15]), 
      .carry(carry[15]));
   FA__1_2550 genblk1_16_F (.a(), .b(y[16]), .cin(carry[15]), .sum(z[16]), 
      .carry(carry[16]));
   FA__1_2547 genblk1_17_F (.a(), .b(y[17]), .cin(carry[16]), .sum(z[17]), 
      .carry(carry[17]));
   FA__1_2544 genblk1_18_F (.a(), .b(y[18]), .cin(carry[17]), .sum(z[18]), 
      .carry(carry[18]));
   FA__1_2541 genblk1_19_F (.a(), .b(y[19]), .cin(carry[18]), .sum(z[19]), 
      .carry(carry[19]));
   FA__1_2538 genblk1_20_F (.a(), .b(y[20]), .cin(carry[19]), .sum(z[20]), 
      .carry(carry[20]));
   FA__1_2535 genblk1_21_F (.a(), .b(y[21]), .cin(carry[20]), .sum(z[21]), 
      .carry(carry[21]));
   FA__1_2532 genblk1_22_F (.a(), .b(y[22]), .cin(carry[21]), .sum(z[22]), 
      .carry(carry[22]));
   FA__1_2529 genblk1_23_F (.a(), .b(y[23]), .cin(carry[22]), .sum(z[23]), 
      .carry(z[24]));
endmodule

module FA__1_881(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_878(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_875(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_872(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_869(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_866(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_863(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_860(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_857(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_854(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_851(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_848(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_845(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_842(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_839(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_836(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_833(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_830(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_827(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_824(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_821(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_815(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_812(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_809(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_806(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_803(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_800(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_797(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_791(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_788(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_785(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_782(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_779(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_776(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_773(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_767(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_764(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_761(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_758(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_755(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_752(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_749(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_743(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_740(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_737(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_734(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_731(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_728(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_725(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_719(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_716(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_713(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_710(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_707(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_704(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_701(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_698(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_695(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_882(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_881 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_878 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_875 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_872 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_869 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_866 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_863 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_860 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_857 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_854 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_851 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_848 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_845 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_842 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_839 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_836 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_833 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_830 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_827 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_824 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_821 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_818 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_815 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_812 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_809 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_806 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_803 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_800 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_797 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_794 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_791 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_788 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_785 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_782 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_779 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_776 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_773 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_770 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_767 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_764 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_761 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_758 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_755 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_752 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_749 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_746 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_743 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_740 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_737 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_734 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_731 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_728 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_725 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_722 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_719 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_716 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_713 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_710 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_707 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_704 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_701 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_698 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_695 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_1135(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1132(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1129(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1126(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1123(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1120(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1117(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1111(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1108(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1105(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1102(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1099(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1096(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1093(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1090(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1087(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1084(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1081(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1078(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1075(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1072(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1069(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1066(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1063(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1060(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1057(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1054(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1051(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1048(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1045(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1042(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1039(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1036(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1033(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1030(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1027(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1024(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1021(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1015(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1012(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1009(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1006(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1003(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1000(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_997(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_991(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_988(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_985(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_982(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_979(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_976(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_973(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_970(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_967(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_964(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_961(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_958(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_955(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_952(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_949(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_1136(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_1135 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_1132 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_1129 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_1126 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_1123 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_1120 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_1117 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_1114 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_1111 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_1108 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_1105 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_1102 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_1099 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_1096 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_1093 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_1090 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_1087 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_1084 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_1081 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_1078 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_1075 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_1072 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_1069 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_1066 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_1063 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_1060 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_1057 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_1054 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_1051 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_1048 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_1045 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_1042 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_1039 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_1036 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_1033 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_1030 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_1027 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_1024 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_1021 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_1018 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_1015 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_1012 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_1009 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_1006 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_1003 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_1000 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_997 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_994 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_991 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_988 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_985 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_982 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_979 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_976 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_973 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_970 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_967 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_964 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_961 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_958 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_955 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_952 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_949 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_2719(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_2716(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2713(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2710(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2707(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2704(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2701(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2695(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2692(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2689(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2686(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2683(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2680(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2677(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2674(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_2792(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_2719 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(), .sum(z[24]), .carry(
      carry[24]));
   FA__1_2716 genblk1_25_F (.a(x[25]), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__1_2713 genblk1_26_F (.a(x[26]), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__1_2710 genblk1_27_F (.a(x[27]), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__1_2707 genblk1_28_F (.a(x[28]), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__1_2704 genblk1_29_F (.a(x[29]), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__1_2701 genblk1_30_F (.a(x[30]), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__1_2698 genblk1_31_F (.a(x[31]), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__1_2695 genblk1_32_F (.a(), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__1_2692 genblk1_33_F (.a(), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__1_2689 genblk1_34_F (.a(), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__1_2686 genblk1_35_F (.a(), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__1_2683 genblk1_36_F (.a(), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__1_2680 genblk1_37_F (.a(), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__1_2677 genblk1_38_F (.a(), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__1_2674 genblk1_39_F (.a(), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(z[40]));
endmodule

module FA__1_2936(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_2933(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2930(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2927(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2924(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2921(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2918(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2915(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2912(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2909(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2906(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2903(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2900(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2897(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2894(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2891(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2888(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2885(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2882(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2879(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2876(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2873(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2870(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2867(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_2864(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_2985(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_2936 genblk1_16_F (.a(x[16]), .b(y[16]), .cin(), .sum(z[16]), .carry(
      carry[16]));
   FA__1_2933 genblk1_17_F (.a(x[17]), .b(y[17]), .cin(carry[16]), .sum(z[17]), 
      .carry(carry[17]));
   FA__1_2930 genblk1_18_F (.a(x[18]), .b(y[18]), .cin(carry[17]), .sum(z[18]), 
      .carry(carry[18]));
   FA__1_2927 genblk1_19_F (.a(x[19]), .b(y[19]), .cin(carry[18]), .sum(z[19]), 
      .carry(carry[19]));
   FA__1_2924 genblk1_20_F (.a(x[20]), .b(y[20]), .cin(carry[19]), .sum(z[20]), 
      .carry(carry[20]));
   FA__1_2921 genblk1_21_F (.a(x[21]), .b(y[21]), .cin(carry[20]), .sum(z[21]), 
      .carry(carry[21]));
   FA__1_2918 genblk1_22_F (.a(x[22]), .b(y[22]), .cin(carry[21]), .sum(z[22]), 
      .carry(carry[22]));
   FA__1_2915 genblk1_23_F (.a(x[23]), .b(y[23]), .cin(carry[22]), .sum(z[23]), 
      .carry(carry[23]));
   FA__1_2912 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(carry[23]), .sum(z[24]), 
      .carry(carry[24]));
   FA__1_2909 genblk1_25_F (.a(), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__1_2906 genblk1_26_F (.a(), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__1_2903 genblk1_27_F (.a(), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__1_2900 genblk1_28_F (.a(), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__1_2897 genblk1_29_F (.a(), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__1_2894 genblk1_30_F (.a(), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__1_2891 genblk1_31_F (.a(), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__1_2888 genblk1_32_F (.a(), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__1_2885 genblk1_33_F (.a(), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__1_2882 genblk1_34_F (.a(), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__1_2879 genblk1_35_F (.a(), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__1_2876 genblk1_36_F (.a(), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__1_2873 genblk1_37_F (.a(), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__1_2870 genblk1_38_F (.a(), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__1_2867 genblk1_39_F (.a(), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__1_2864 genblk1_40_F (.a(), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(z[41]));
endmodule

module FA__1_1389(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1383(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1380(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1377(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1374(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1371(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1368(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1365(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1359(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1356(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1353(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1350(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1347(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1344(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1341(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1335(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1332(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1329(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1326(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1323(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1320(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1317(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1311(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1308(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1305(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1302(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1299(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1296(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1293(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1287(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1284(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1281(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1278(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1275(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1272(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1269(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1263(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1260(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1257(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1254(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1251(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1248(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1245(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1242(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1239(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1236(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1233(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1230(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1227(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1224(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1221(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1215(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1212(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1209(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1206(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1203(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_1390(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_1389 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_1386 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_1383 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_1380 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_1377 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_1374 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_1371 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_1368 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_1365 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_1362 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_1359 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_1356 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_1353 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_1350 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_1347 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_1344 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_1341 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_1338 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_1335 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_1332 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_1329 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_1326 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_1323 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_1320 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_1317 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_1314 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_1311 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_1308 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_1305 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_1302 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_1299 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_1296 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_1293 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_1290 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_1287 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_1284 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_1281 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_1278 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_1275 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_1272 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_1269 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_1266 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_1263 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_1260 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_1257 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_1254 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_1251 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_1248 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_1245 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_1242 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_1239 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_1236 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_1233 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_1230 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_1227 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_1224 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_1221 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_1218 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_1215 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_1212 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_1209 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_1206 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_1203 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_1643(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1640(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1637(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1634(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1631(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1628(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1625(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1622(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1619(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1616(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1613(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1610(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1607(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1604(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1601(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1598(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1595(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1592(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1589(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1586(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1583(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1580(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1577(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1574(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1571(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1568(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1565(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1559(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1556(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1553(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1550(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1547(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1544(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1541(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1538(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1535(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1532(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1529(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1526(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1523(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1520(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1517(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1511(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1508(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1505(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1502(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1499(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1496(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1493(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1490(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1487(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1484(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1481(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1478(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1475(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1472(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1469(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1463(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1460(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1457(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_1644(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_1643 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_1640 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_1637 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_1634 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_1631 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_1628 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_1625 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_1622 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_1619 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_1616 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_1613 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_1610 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_1607 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_1604 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_1601 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_1598 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_1595 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_1592 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_1589 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_1586 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_1583 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_1580 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_1577 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_1574 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_1571 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_1568 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_1565 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_1562 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_1559 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_1556 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_1553 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_1550 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_1547 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_1544 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_1541 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_1538 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_1535 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_1532 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_1529 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_1526 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_1523 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_1520 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_1517 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_1514 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_1511 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_1508 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_1505 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_1502 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_1499 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_1496 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_1493 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_1490 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_1487 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_1484 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_1481 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_1478 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_1475 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_1472 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_1469 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_1466 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_1463 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_1460 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_1457 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_3129(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_3126(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3123(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3120(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3117(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3111(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3108(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3105(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3102(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3099(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3096(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3093(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3090(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3087(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3084(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_3178(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_3129 genblk1_16_F (.a(x[16]), .b(y[16]), .cin(), .sum(z[16]), .carry(
      carry[16]));
   FA__1_3126 genblk1_17_F (.a(x[17]), .b(y[17]), .cin(carry[16]), .sum(z[17]), 
      .carry(carry[17]));
   FA__1_3123 genblk1_18_F (.a(x[18]), .b(y[18]), .cin(carry[17]), .sum(z[18]), 
      .carry(carry[18]));
   FA__1_3120 genblk1_19_F (.a(x[19]), .b(y[19]), .cin(carry[18]), .sum(z[19]), 
      .carry(carry[19]));
   FA__1_3117 genblk1_20_F (.a(x[20]), .b(y[20]), .cin(carry[19]), .sum(z[20]), 
      .carry(carry[20]));
   FA__1_3114 genblk1_21_F (.a(x[21]), .b(y[21]), .cin(carry[20]), .sum(z[21]), 
      .carry(carry[21]));
   FA__1_3111 genblk1_22_F (.a(x[22]), .b(y[22]), .cin(carry[21]), .sum(z[22]), 
      .carry(carry[22]));
   FA__1_3108 genblk1_23_F (.a(x[23]), .b(y[23]), .cin(carry[22]), .sum(z[23]), 
      .carry(carry[23]));
   FA__1_3105 genblk1_24_F (.a(), .b(y[24]), .cin(carry[23]), .sum(z[24]), 
      .carry(carry[24]));
   FA__1_3102 genblk1_25_F (.a(), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__1_3099 genblk1_26_F (.a(), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__1_3096 genblk1_27_F (.a(), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__1_3093 genblk1_28_F (.a(), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__1_3090 genblk1_29_F (.a(), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__1_3087 genblk1_30_F (.a(), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__1_3084 genblk1_31_F (.a(), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(z[32]));
endmodule

module FA__1_1897(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1894(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1891(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1888(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1885(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1882(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1879(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1876(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1873(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1870(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1867(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1864(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1861(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1858(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1855(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1852(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_1849(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1846(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1843(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1840(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1837(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1831(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1828(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1825(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1822(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1819(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1816(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1813(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1807(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1804(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1801(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1798(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1795(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1792(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1789(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1783(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1780(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1777(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1774(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1771(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1768(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1765(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1759(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1756(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1753(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1750(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1747(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1744(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1741(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1735(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1732(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1729(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1726(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1723(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1720(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1717(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1714(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1711(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_1898(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_1897 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_1894 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_1891 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_1888 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_1885 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_1882 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_1879 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_1876 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_1873 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_1870 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_1867 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_1864 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_1861 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_1858 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_1855 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_1852 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_1849 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_1846 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_1843 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_1840 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_1837 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_1834 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_1831 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_1828 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_1825 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_1822 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_1819 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_1816 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_1813 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_1810 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_1807 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_1804 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_1801 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_1798 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_1795 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_1792 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_1789 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_1786 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_1783 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_1780 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_1777 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_1774 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_1771 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_1768 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_1765 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_1762 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_1759 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_1756 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_1753 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_1750 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_1747 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_1744 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_1741 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_1738 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_1735 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_1732 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_1729 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_1726 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_1723 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_1720 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_1717 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_1714 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_1711 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_2151(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2148(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2145(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2142(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2139(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2136(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2133(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2127(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2124(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2121(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2118(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2115(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2112(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2109(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2106(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2103(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2100(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2097(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2094(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2091(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2088(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2085(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2082(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2079(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2076(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2073(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2070(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2067(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2064(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2061(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2058(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2055(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2052(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2049(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2046(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2043(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2040(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2037(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2034(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2031(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2028(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2025(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2022(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2019(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2016(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2013(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2010(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2007(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2004(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2001(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1998(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1995(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1992(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1989(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1986(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1983(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1980(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1977(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1974(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_1971(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_1968(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_1965(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_2152(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_2151 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_2148 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_2145 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_2142 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_2139 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_2136 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_2133 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_2130 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_2127 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_2124 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_2121 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_2118 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_2115 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_2112 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_2109 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_2106 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_2103 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_2100 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_2097 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_2094 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_2091 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_2088 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_2085 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_2082 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_2079 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_2076 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_2073 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_2070 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_2067 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_2064 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_2061 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_2058 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_2055 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_2052 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_2049 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_2046 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_2043 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_2040 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_2037 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_2034 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_2031 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_2028 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_2025 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_2022 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_2019 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_2016 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_2013 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_2010 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_2007 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_2004 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_2001 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_1998 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_1995 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_1992 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_1989 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_1986 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_1983 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_1980 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_1977 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_1974 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_1971 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_1968 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_1965 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__1_3274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_3271(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3268(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3265(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3262(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3259(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3256(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3253(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3247(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3244(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3241(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3238(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3235(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3232(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3229(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_3371(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_3274 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(), .sum(z[32]), .carry(
      carry[32]));
   FA__1_3271 genblk1_33_F (.a(x[33]), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__1_3268 genblk1_34_F (.a(x[34]), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__1_3265 genblk1_35_F (.a(x[35]), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__1_3262 genblk1_36_F (.a(x[36]), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__1_3259 genblk1_37_F (.a(x[37]), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__1_3256 genblk1_38_F (.a(x[38]), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__1_3253 genblk1_39_F (.a(x[39]), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__1_3250 genblk1_40_F (.a(), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__1_3247 genblk1_41_F (.a(), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__1_3244 genblk1_42_F (.a(), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__1_3241 genblk1_43_F (.a(), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__1_3238 genblk1_44_F (.a(), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__1_3235 genblk1_45_F (.a(), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__1_3232 genblk1_46_F (.a(), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__1_3229 genblk1_47_F (.a(), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(z[48]));
endmodule

module FA__1_3491(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_3488(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3485(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3482(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3479(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3476(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3473(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3470(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3467(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3464(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3461(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3458(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3455(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3452(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3449(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3446(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3443(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3440(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3437(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3434(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3431(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3428(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3425(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3422(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3419(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_3564(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_3491 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(), .sum(z[24]), .carry(
      carry[24]));
   FA__1_3488 genblk1_25_F (.a(x[25]), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__1_3485 genblk1_26_F (.a(x[26]), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__1_3482 genblk1_27_F (.a(x[27]), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__1_3479 genblk1_28_F (.a(x[28]), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__1_3476 genblk1_29_F (.a(x[29]), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__1_3473 genblk1_30_F (.a(x[30]), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__1_3470 genblk1_31_F (.a(x[31]), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__1_3467 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__1_3464 genblk1_33_F (.a(), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__1_3461 genblk1_34_F (.a(), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__1_3458 genblk1_35_F (.a(), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__1_3455 genblk1_36_F (.a(), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__1_3452 genblk1_37_F (.a(), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__1_3449 genblk1_38_F (.a(), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__1_3446 genblk1_39_F (.a(), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__1_3443 genblk1_40_F (.a(), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__1_3440 genblk1_41_F (.a(), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__1_3437 genblk1_42_F (.a(), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__1_3434 genblk1_43_F (.a(), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__1_3431 genblk1_44_F (.a(), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__1_3428 genblk1_45_F (.a(), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__1_3425 genblk1_46_F (.a(), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__1_3422 genblk1_47_F (.a(), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__1_3419 genblk1_48_F (.a(), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(z[49]));
endmodule

module FA__1_3732(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_3729(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3726(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3723(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3720(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3717(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3711(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3708(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3705(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3702(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3699(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3696(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3693(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3690(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3687(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3684(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3681(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3678(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3675(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3672(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3669(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3666(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3663(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3660(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3657(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3654(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3651(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3648(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3645(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3642(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3639(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3636(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3633(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_3630(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3627(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3624(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3621(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3615(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3612(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_3609(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__1_3757(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_3732 genblk1_8_F (.a(x[8]), .b(y[8]), .cin(), .sum(z[8]), .carry(
      carry[8]));
   FA__1_3729 genblk1_9_F (.a(x[9]), .b(y[9]), .cin(carry[8]), .sum(z[9]), 
      .carry(carry[9]));
   FA__1_3726 genblk1_10_F (.a(x[10]), .b(y[10]), .cin(carry[9]), .sum(z[10]), 
      .carry(carry[10]));
   FA__1_3723 genblk1_11_F (.a(x[11]), .b(y[11]), .cin(carry[10]), .sum(z[11]), 
      .carry(carry[11]));
   FA__1_3720 genblk1_12_F (.a(x[12]), .b(y[12]), .cin(carry[11]), .sum(z[12]), 
      .carry(carry[12]));
   FA__1_3717 genblk1_13_F (.a(x[13]), .b(y[13]), .cin(carry[12]), .sum(z[13]), 
      .carry(carry[13]));
   FA__1_3714 genblk1_14_F (.a(x[14]), .b(y[14]), .cin(carry[13]), .sum(z[14]), 
      .carry(carry[14]));
   FA__1_3711 genblk1_15_F (.a(x[15]), .b(y[15]), .cin(carry[14]), .sum(z[15]), 
      .carry(carry[15]));
   FA__1_3708 genblk1_16_F (.a(x[16]), .b(y[16]), .cin(carry[15]), .sum(z[16]), 
      .carry(carry[16]));
   FA__1_3705 genblk1_17_F (.a(x[17]), .b(y[17]), .cin(carry[16]), .sum(z[17]), 
      .carry(carry[17]));
   FA__1_3702 genblk1_18_F (.a(x[18]), .b(y[18]), .cin(carry[17]), .sum(z[18]), 
      .carry(carry[18]));
   FA__1_3699 genblk1_19_F (.a(x[19]), .b(y[19]), .cin(carry[18]), .sum(z[19]), 
      .carry(carry[19]));
   FA__1_3696 genblk1_20_F (.a(x[20]), .b(y[20]), .cin(carry[19]), .sum(z[20]), 
      .carry(carry[20]));
   FA__1_3693 genblk1_21_F (.a(x[21]), .b(y[21]), .cin(carry[20]), .sum(z[21]), 
      .carry(carry[21]));
   FA__1_3690 genblk1_22_F (.a(x[22]), .b(y[22]), .cin(carry[21]), .sum(z[22]), 
      .carry(carry[22]));
   FA__1_3687 genblk1_23_F (.a(x[23]), .b(y[23]), .cin(carry[22]), .sum(z[23]), 
      .carry(carry[23]));
   FA__1_3684 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(carry[23]), .sum(z[24]), 
      .carry(carry[24]));
   FA__1_3681 genblk1_25_F (.a(x[25]), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__1_3678 genblk1_26_F (.a(x[26]), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__1_3675 genblk1_27_F (.a(x[27]), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__1_3672 genblk1_28_F (.a(x[28]), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__1_3669 genblk1_29_F (.a(x[29]), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__1_3666 genblk1_30_F (.a(x[30]), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__1_3663 genblk1_31_F (.a(x[31]), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__1_3660 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__1_3657 genblk1_33_F (.a(x[33]), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__1_3654 genblk1_34_F (.a(x[34]), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__1_3651 genblk1_35_F (.a(x[35]), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__1_3648 genblk1_36_F (.a(x[36]), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__1_3645 genblk1_37_F (.a(x[37]), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__1_3642 genblk1_38_F (.a(x[38]), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__1_3639 genblk1_39_F (.a(x[39]), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__1_3636 genblk1_40_F (.a(x[40]), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__1_3633 genblk1_41_F (.a(x[41]), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__1_3630 genblk1_42_F (.a(), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__1_3627 genblk1_43_F (.a(), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__1_3624 genblk1_44_F (.a(), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__1_3621 genblk1_45_F (.a(), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__1_3618 genblk1_46_F (.a(), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__1_3615 genblk1_47_F (.a(), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__1_3612 genblk1_48_F (.a(), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(carry[48]));
   FA__1_3609 genblk1_49_F (.a(), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(z[50]));
endmodule

module datapath__0_81(p_0, B);
   output [31:0]p_0;
   input [31:0]B;

   XOR2_X1 i_0 (.A(B[1]), .B(B[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(B[2]), .B1(B[1]), .B2(B[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(B[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(B[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(B[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(B[6]), .B1(n_27), .B2(B[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(B[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(B[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(B[9]), .B1(n_25), .B2(B[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(B[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(B[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(B[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(B[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(B[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(B[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(B[16]), .B1(n_19), .B2(B[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(B[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(B[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(B[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(B[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(B[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(B[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(B[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(B[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(B[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(B[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(B[27]), .B1(n_9), .B2(B[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(B[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(B[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(B[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(B[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(B[28]), .A3(B[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(B[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(B[26]), .A3(B[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(B[23]), .A3(B[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(B[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(B[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(B[18]), .A3(B[19]), .A4(B[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(B[18]), .A3(B[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(B[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(B[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(B[15]), .A3(B[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(B[12]), .A3(B[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(B[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(B[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(B[8]), .A3(B[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(B[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(B[5]), .A3(B[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(B[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(B[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(B[2]), .A2(B[1]), .A3(B[0]), .ZN(n_29));
   INV_X1 i_61 (.A(B[11]), .ZN(n_30));
   INV_X1 i_62 (.A(B[14]), .ZN(n_31));
   INV_X1 i_63 (.A(B[21]), .ZN(n_32));
   INV_X1 i_64 (.A(B[25]), .ZN(n_33));
endmodule

module datapath__0_79(p_0, A);
   output [31:0]p_0;
   input [31:0]A;

   XOR2_X1 i_0 (.A(A[1]), .B(A[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(A[2]), .B1(A[1]), .B2(A[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(A[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(A[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(A[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(A[6]), .B1(n_27), .B2(A[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(A[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(A[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(A[9]), .B1(n_25), .B2(A[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(A[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(A[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(A[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(A[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(A[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(A[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(A[16]), .B1(n_19), .B2(A[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(A[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(A[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(A[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(A[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(A[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(A[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(A[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(A[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(A[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(A[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(A[27]), .B1(n_9), .B2(A[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(A[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(A[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(A[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(A[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(A[28]), .A3(A[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(A[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(A[26]), .A3(A[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(A[23]), .A3(A[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(A[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(A[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(A[18]), .A3(A[19]), .A4(A[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(A[18]), .A3(A[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(A[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(A[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(A[15]), .A3(A[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(A[12]), .A3(A[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(A[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(A[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(A[8]), .A3(A[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(A[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(A[5]), .A3(A[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(A[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(A[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(A[2]), .A2(A[1]), .A3(A[0]), .ZN(n_29));
   INV_X1 i_61 (.A(A[11]), .ZN(n_30));
   INV_X1 i_62 (.A(A[14]), .ZN(n_31));
   INV_X1 i_63 (.A(A[21]), .ZN(n_32));
   INV_X1 i_64 (.A(A[25]), .ZN(n_33));
endmodule

module FA__1_2405(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2402(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2399(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2396(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2393(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2390(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2387(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2384(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2381(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2378(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2375(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2372(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2369(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2366(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2363(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2360(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_2357(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2351(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2348(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2345(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2342(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2339(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2336(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2333(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2327(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2324(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2321(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2318(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2315(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2312(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2309(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2303(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2300(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2297(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2294(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2291(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2288(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2285(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2279(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2276(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2273(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2270(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2267(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2264(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2261(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2258(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2255(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2252(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2249(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2246(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2243(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2240(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2237(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2231(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2228(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_2225(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_2222(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_2219(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__1_2406(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_2405 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_2402 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_2399 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_2396 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_2393 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_2390 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_2387 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_2384 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_2381 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_2378 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_2375 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_2372 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_2369 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_2366 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_2363 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_2360 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_2357 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_2354 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_2351 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_2348 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_2345 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_2342 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_2339 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_2336 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_2333 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_2330 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_2327 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_2324 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_2321 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_2318 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_2315 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_2312 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_2309 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_2306 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_2303 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_2300 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_2297 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_2294 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_2291 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_2288 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_2285 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_2282 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_2279 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_2276 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_2273 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_2270 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_2267 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_2264 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_2261 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_2258 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_2255 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_2252 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_2249 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_2246 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_2243 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_2240 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_2237 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_2234 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_2231 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_2228 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_2225 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_2222 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_2219 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module datapath(p_0, out);
   output [63:0]p_0;
   input [63:0]out;

   XOR2_X1 i_0 (.A(out[1]), .B(out[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(out[2]), .B1(out[1]), .B2(out[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(out[3]), .B(n_61), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(out[4]), .B(n_60), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(out[5]), .B(n_59), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(out[6]), .B1(n_59), .B2(out[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(out[7]), .B(n_58), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(out[8]), .B(n_57), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(out[9]), .B1(n_57), .B2(out[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(out[10]), .B(n_56), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(out[11]), .B(n_55), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(out[12]), .B(n_54), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(out[13]), .B(n_53), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(out[14]), .B(n_52), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(out[15]), .B1(n_52), .B2(out[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(out[16]), .B(n_51), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(out[17]), .B(n_50), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(out[18]), .B(n_49), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(out[19]), .B(n_48), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(out[20]), .B(n_47), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(out[21]), .B(n_46), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(out[22]), .B(n_45), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(out[23]), .B(n_44), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(out[24]), .B(n_43), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(out[25]), .B(n_42), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(out[26]), .B(n_41), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(out[27]), .B(n_40), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(out[28]), .B(n_39), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(out[29]), .B(n_38), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(out[30]), .B(n_37), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(out[31]), .B(n_36), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(out[32]), .B(n_35), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(out[33]), .B(n_34), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(out[34]), .B(n_33), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(out[35]), .B(n_32), .ZN(p_0[35]));
   XNOR2_X1 i_39 (.A(out[36]), .B(n_31), .ZN(p_0[36]));
   XOR2_X1 i_40 (.A(out[37]), .B(n_30), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(out[38]), .B(n_29), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(out[39]), .B(n_28), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(out[40]), .B(n_27), .ZN(p_0[40]));
   XOR2_X1 i_44 (.A(out[41]), .B(n_26), .Z(p_0[41]));
   XNOR2_X1 i_45 (.A(out[42]), .B(n_25), .ZN(p_0[42]));
   XOR2_X1 i_46 (.A(out[43]), .B(n_24), .Z(p_0[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(p_0[44]));
   OAI21_X1 i_48 (.A(out[44]), .B1(n_24), .B2(out[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(out[45]), .B(n_23), .Z(p_0[45]));
   XOR2_X1 i_50 (.A(out[46]), .B(n_22), .Z(p_0[46]));
   XOR2_X1 i_51 (.A(out[47]), .B(n_21), .Z(p_0[47]));
   XOR2_X1 i_52 (.A(out[48]), .B(n_20), .Z(p_0[48]));
   XNOR2_X1 i_53 (.A(out[49]), .B(n_19), .ZN(p_0[49]));
   XNOR2_X1 i_54 (.A(out[50]), .B(n_18), .ZN(p_0[50]));
   XNOR2_X1 i_55 (.A(out[51]), .B(n_17), .ZN(p_0[51]));
   XOR2_X1 i_56 (.A(out[52]), .B(n_16), .Z(p_0[52]));
   XNOR2_X1 i_57 (.A(out[53]), .B(n_15), .ZN(p_0[53]));
   XNOR2_X1 i_58 (.A(out[54]), .B(n_14), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(out[55]), .B(n_13), .ZN(p_0[55]));
   XOR2_X1 i_60 (.A(out[56]), .B(n_12), .Z(p_0[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(p_0[57]));
   OAI21_X1 i_62 (.A(out[57]), .B1(n_12), .B2(out[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(out[58]), .B(n_11), .Z(p_0[58]));
   XNOR2_X1 i_64 (.A(out[59]), .B(n_10), .ZN(p_0[59]));
   XNOR2_X1 i_65 (.A(out[60]), .B(n_9), .ZN(p_0[60]));
   XOR2_X1 i_66 (.A(out[61]), .B(n_8), .Z(p_0[61]));
   XNOR2_X1 i_67 (.A(out[62]), .B(n_7), .ZN(p_0[62]));
   XNOR2_X1 i_68 (.A(out[63]), .B(n_6), .ZN(p_0[63]));
   NOR3_X1 i_69 (.A1(n_8), .A2(out[61]), .A3(out[62]), .ZN(n_6));
   NOR2_X1 i_70 (.A1(n_8), .A2(out[61]), .ZN(n_7));
   NAND2_X1 i_71 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_72 (.A1(n_11), .A2(out[58]), .A3(out[59]), .ZN(n_9));
   NOR2_X1 i_73 (.A1(n_11), .A2(out[58]), .ZN(n_10));
   OR3_X1 i_74 (.A1(n_12), .A2(out[56]), .A3(out[57]), .ZN(n_11));
   NAND2_X1 i_75 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_76 (.A1(n_16), .A2(out[52]), .A3(out[53]), .A4(out[54]), .ZN(n_13));
   NOR3_X1 i_77 (.A1(n_16), .A2(out[52]), .A3(out[53]), .ZN(n_14));
   NOR2_X1 i_78 (.A1(n_16), .A2(out[52]), .ZN(n_15));
   NAND2_X1 i_79 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_80 (.A1(n_20), .A2(out[48]), .A3(out[49]), .A4(out[50]), .ZN(n_17));
   NOR3_X1 i_81 (.A1(n_20), .A2(out[48]), .A3(out[49]), .ZN(n_18));
   NOR2_X1 i_82 (.A1(n_20), .A2(out[48]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(out[47]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(out[46]), .ZN(n_21));
   OR2_X1 i_85 (.A1(n_23), .A2(out[45]), .ZN(n_22));
   OR3_X1 i_86 (.A1(n_24), .A2(out[43]), .A3(out[44]), .ZN(n_23));
   NAND2_X1 i_87 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_88 (.A1(n_26), .A2(out[41]), .ZN(n_25));
   NAND2_X1 i_89 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_90 (.A1(n_29), .A2(out[38]), .A3(out[39]), .ZN(n_27));
   NOR2_X1 i_91 (.A1(n_29), .A2(out[38]), .ZN(n_28));
   OR2_X1 i_92 (.A1(n_30), .A2(out[37]), .ZN(n_29));
   NAND2_X1 i_93 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_94 (.A1(n_34), .A2(out[33]), .A3(out[34]), .A4(out[35]), .ZN(n_31));
   NOR3_X1 i_95 (.A1(n_34), .A2(out[33]), .A3(out[34]), .ZN(n_32));
   NOR2_X1 i_96 (.A1(n_34), .A2(out[33]), .ZN(n_33));
   OR2_X1 i_97 (.A1(n_35), .A2(out[32]), .ZN(n_34));
   NAND2_X1 i_98 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_99 (.A1(n_39), .A2(out[28]), .A3(out[29]), .A4(out[30]), .ZN(n_36));
   NOR3_X1 i_100 (.A1(n_39), .A2(out[28]), .A3(out[29]), .ZN(n_37));
   NOR2_X1 i_101 (.A1(n_39), .A2(out[28]), .ZN(n_38));
   OR2_X1 i_102 (.A1(n_40), .A2(out[27]), .ZN(n_39));
   NAND2_X1 i_103 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_104 (.A1(n_44), .A2(out[23]), .A3(out[24]), .A4(out[25]), .ZN(n_41));
   NOR3_X1 i_105 (.A1(n_44), .A2(out[23]), .A3(out[24]), .ZN(n_42));
   NOR2_X1 i_106 (.A1(n_44), .A2(out[23]), .ZN(n_43));
   OR2_X1 i_107 (.A1(n_45), .A2(out[22]), .ZN(n_44));
   NAND2_X1 i_108 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_109 (.A1(n_49), .A2(out[18]), .A3(out[19]), .A4(out[20]), .ZN(n_46));
   NOR3_X1 i_110 (.A1(n_49), .A2(out[18]), .A3(out[19]), .ZN(n_47));
   NOR2_X1 i_111 (.A1(n_49), .A2(out[18]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(out[17]), .ZN(n_49));
   OR2_X1 i_113 (.A1(n_51), .A2(out[16]), .ZN(n_50));
   OR3_X1 i_114 (.A1(n_52), .A2(out[14]), .A3(out[15]), .ZN(n_51));
   NAND2_X1 i_115 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_116 (.A1(n_54), .A2(out[12]), .ZN(n_53));
   NAND2_X1 i_117 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_118 (.A1(n_56), .A2(out[10]), .ZN(n_55));
   OR3_X1 i_119 (.A1(n_57), .A2(out[8]), .A3(out[9]), .ZN(n_56));
   OR2_X1 i_120 (.A1(n_58), .A2(out[7]), .ZN(n_57));
   OR3_X1 i_121 (.A1(n_59), .A2(out[5]), .A3(out[6]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(out[4]), .ZN(n_59));
   OR2_X1 i_123 (.A1(n_61), .A2(out[3]), .ZN(n_60));
   OR3_X1 i_124 (.A1(out[2]), .A2(out[1]), .A3(out[0]), .ZN(n_61));
   INV_X1 i_125 (.A(out[11]), .ZN(n_62));
   INV_X1 i_126 (.A(out[13]), .ZN(n_63));
   INV_X1 i_127 (.A(out[21]), .ZN(n_64));
   INV_X1 i_128 (.A(out[26]), .ZN(n_65));
   INV_X1 i_129 (.A(out[31]), .ZN(n_66));
   INV_X1 i_130 (.A(out[36]), .ZN(n_67));
   INV_X1 i_131 (.A(out[40]), .ZN(n_68));
   INV_X1 i_132 (.A(out[42]), .ZN(n_69));
   INV_X1 i_133 (.A(out[51]), .ZN(n_70));
   INV_X1 i_134 (.A(out[55]), .ZN(n_71));
   INV_X1 i_135 (.A(out[60]), .ZN(n_72));
endmodule

module FA__1_188(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__1_191(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_197(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_200(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_203(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_206(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_209(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_212(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_215(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_221(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_224(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_227(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_230(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_233(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_236(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_239(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_245(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_248(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_251(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_254(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_257(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_260(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_263(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_269(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_272(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_275(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_278(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_281(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_284(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_287(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_293(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_296(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_299(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_302(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_305(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_308(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_311(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_317(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_320(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_323(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__1_326(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__0_149(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(sum));
endmodule

module adder64__0_154(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__1_188 genblk1_16_F (.a(x[16]), .b(y[16]), .cin(), .sum(z[16]), .carry(
      carry[16]));
   FA__1_191 genblk1_17_F (.a(x[17]), .b(y[17]), .cin(carry[16]), .sum(z[17]), 
      .carry(carry[17]));
   FA__1_194 genblk1_18_F (.a(x[18]), .b(y[18]), .cin(carry[17]), .sum(z[18]), 
      .carry(carry[18]));
   FA__1_197 genblk1_19_F (.a(x[19]), .b(y[19]), .cin(carry[18]), .sum(z[19]), 
      .carry(carry[19]));
   FA__1_200 genblk1_20_F (.a(x[20]), .b(y[20]), .cin(carry[19]), .sum(z[20]), 
      .carry(carry[20]));
   FA__1_203 genblk1_21_F (.a(x[21]), .b(y[21]), .cin(carry[20]), .sum(z[21]), 
      .carry(carry[21]));
   FA__1_206 genblk1_22_F (.a(x[22]), .b(y[22]), .cin(carry[21]), .sum(z[22]), 
      .carry(carry[22]));
   FA__1_209 genblk1_23_F (.a(x[23]), .b(y[23]), .cin(carry[22]), .sum(z[23]), 
      .carry(carry[23]));
   FA__1_212 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(carry[23]), .sum(z[24]), 
      .carry(carry[24]));
   FA__1_215 genblk1_25_F (.a(x[25]), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__1_218 genblk1_26_F (.a(x[26]), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__1_221 genblk1_27_F (.a(x[27]), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__1_224 genblk1_28_F (.a(x[28]), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__1_227 genblk1_29_F (.a(x[29]), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__1_230 genblk1_30_F (.a(x[30]), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__1_233 genblk1_31_F (.a(x[31]), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__1_236 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__1_239 genblk1_33_F (.a(x[33]), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__1_242 genblk1_34_F (.a(x[34]), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__1_245 genblk1_35_F (.a(x[35]), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__1_248 genblk1_36_F (.a(x[36]), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__1_251 genblk1_37_F (.a(x[37]), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__1_254 genblk1_38_F (.a(x[38]), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__1_257 genblk1_39_F (.a(x[39]), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__1_260 genblk1_40_F (.a(x[40]), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__1_263 genblk1_41_F (.a(x[41]), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__1_266 genblk1_42_F (.a(x[42]), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__1_269 genblk1_43_F (.a(x[43]), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__1_272 genblk1_44_F (.a(x[44]), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__1_275 genblk1_45_F (.a(x[45]), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__1_278 genblk1_46_F (.a(x[46]), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__1_281 genblk1_47_F (.a(x[47]), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__1_284 genblk1_48_F (.a(x[48]), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(carry[48]));
   FA__1_287 genblk1_49_F (.a(x[49]), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(carry[49]));
   FA__1_290 genblk1_50_F (.a(x[50]), .b(y[50]), .cin(carry[49]), .sum(z[50]), 
      .carry(carry[50]));
   FA__1_293 genblk1_51_F (.a(), .b(y[51]), .cin(carry[50]), .sum(z[51]), 
      .carry(carry[51]));
   FA__1_296 genblk1_52_F (.a(), .b(y[52]), .cin(carry[51]), .sum(z[52]), 
      .carry(carry[52]));
   FA__1_299 genblk1_53_F (.a(), .b(y[53]), .cin(carry[52]), .sum(z[53]), 
      .carry(carry[53]));
   FA__1_302 genblk1_54_F (.a(), .b(y[54]), .cin(carry[53]), .sum(z[54]), 
      .carry(carry[54]));
   FA__1_305 genblk1_55_F (.a(), .b(y[55]), .cin(carry[54]), .sum(z[55]), 
      .carry(carry[55]));
   FA__1_308 genblk1_56_F (.a(), .b(y[56]), .cin(carry[55]), .sum(z[56]), 
      .carry(carry[56]));
   FA__1_311 genblk1_57_F (.a(), .b(y[57]), .cin(carry[56]), .sum(z[57]), 
      .carry(carry[57]));
   FA__1_314 genblk1_58_F (.a(), .b(y[58]), .cin(carry[57]), .sum(z[58]), 
      .carry(carry[58]));
   FA__1_317 genblk1_59_F (.a(), .b(y[59]), .cin(carry[58]), .sum(z[59]), 
      .carry(carry[59]));
   FA__1_320 genblk1_60_F (.a(), .b(y[60]), .cin(carry[59]), .sum(z[60]), 
      .carry(carry[60]));
   FA__1_323 genblk1_61_F (.a(), .b(y[61]), .cin(carry[60]), .sum(z[61]), 
      .carry(carry[61]));
   FA__1_326 genblk1_62_F (.a(), .b(y[62]), .cin(carry[61]), .sum(z[62]), 
      .carry(carry[62]));
   FA__0_149 genblk1_63_F (.a(), .b(y[63]), .cin(carry[62]), .sum(z[63]), .carry());
endmodule

module FA__1_2(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_5(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_8(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_11(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_14(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_329(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_17(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_20(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_23(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_26(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_332(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_335(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_338(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_341(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_344(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_347(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__1_350(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_29(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_32(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_35(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_353(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_38(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_356(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_41(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_44(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_47(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_50(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_53(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_56(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_59(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_62(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_359(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_65(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_68(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_71(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_74(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_77(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_80(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_83(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_86(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_89(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_92(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_95(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_98(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_101(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_104(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_107(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_110(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_113(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_362(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_116(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_365(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_119(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_122(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_125(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_368(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_128(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_131(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_371(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_134(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__1_137(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__1_374(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__1_140(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__0_153(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__1_2 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__1_5 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__1_8 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__1_11 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__1_14 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__1_329 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__1_17 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__1_20 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__1_23 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__1_26 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__1_332 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__1_335 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__1_338 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__1_341 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__1_344 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__1_347 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__1_350 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__1_29 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__1_32 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__1_35 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__1_353 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__1_38 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__1_356 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__1_41 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__1_44 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__1_47 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__1_50 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__1_53 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__1_56 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__1_59 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__1_62 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__1_359 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__1_65 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__1_68 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__1_71 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__1_74 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__1_77 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__1_80 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__1_83 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__1_86 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__1_89 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__1_92 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__1_95 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__1_98 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__1_101 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__1_104 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__1_107 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__1_110 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__1_113 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__1_362 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__1_116 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__1_365 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__1_119 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__1_122 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__1_125 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__1_368 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__1_128 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__1_131 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__1_371 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__1_134 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__1_137 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__1_374 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__1_140 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_1994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_1991(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1988(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1985(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1982(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1979(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1976(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1973(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1970(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1967(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1964(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1961(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1958(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1955(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1952(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_1949(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__2_2091(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_1994 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(), .sum(z[32]), .carry(
      carry[32]));
   FA__2_1991 genblk1_33_F (.a(x[33]), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__2_1988 genblk1_34_F (.a(x[34]), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__2_1985 genblk1_35_F (.a(x[35]), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__2_1982 genblk1_36_F (.a(x[36]), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__2_1979 genblk1_37_F (.a(x[37]), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__2_1976 genblk1_38_F (.a(x[38]), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__2_1973 genblk1_39_F (.a(x[39]), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__2_1970 genblk1_40_F (.a(), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__2_1967 genblk1_41_F (.a(), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__2_1964 genblk1_42_F (.a(), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__2_1961 genblk1_43_F (.a(), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__2_1958 genblk1_44_F (.a(), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__2_1955 genblk1_45_F (.a(), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__2_1952 genblk1_46_F (.a(), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__2_1949 genblk1_47_F (.a(), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(z[48]));
endmodule

module FA__2_627(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_624(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_621(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_615(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_612(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_609(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_606(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_603(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_600(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_597(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_594(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_591(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_588(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_585(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_582(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_579(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_576(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_573(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_567(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_564(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_561(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_558(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_555(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_552(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_549(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_546(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_543(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_540(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_537(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_534(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_531(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_528(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_525(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_519(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_516(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_513(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_510(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_507(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_504(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_501(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_495(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_492(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_489(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_486(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_483(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_480(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_477(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_474(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_471(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_468(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_465(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_462(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_459(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_456(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_453(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_447(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_444(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_441(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__2_628(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_627 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_624 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_621 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_618 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_615 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_612 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_609 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_606 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_603 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_600 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_597 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_594 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_591 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_588 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_585 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_582 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_579 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_576 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_573 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_570 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_567 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_564 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_561 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_558 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_555 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_552 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_549 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_546 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_543 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_540 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_537 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_534 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_531 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_528 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_525 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_522 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_519 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_516 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_513 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_510 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_507 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_504 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_501 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_498 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_495 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_492 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_489 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_486 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_483 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_480 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_477 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_474 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_471 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_468 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_465 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_462 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_459 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_456 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_453 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_450 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_447 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_444 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_441 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_881(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_878(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_875(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_872(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_869(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_866(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_863(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_860(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_857(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_854(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_851(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_848(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_845(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_842(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_839(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_836(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_833(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_830(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_827(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_824(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_821(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_815(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_812(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_809(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_806(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_803(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_800(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_797(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_791(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_788(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_785(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_782(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_779(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_776(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_773(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_767(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_764(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_761(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_758(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_755(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_752(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_749(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_743(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_740(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_737(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_734(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_731(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_728(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_725(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_719(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_716(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_713(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_710(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_707(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_704(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_701(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_698(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_695(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__2_882(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_881 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_878 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_875 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_872 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_869 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_866 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_863 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_860 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_857 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_854 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_851 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_848 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_845 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_842 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_839 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_836 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_833 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_830 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_827 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_824 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_821 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_818 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_815 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_812 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_809 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_806 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_803 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_800 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_797 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_794 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_791 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_788 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_785 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_782 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_779 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_776 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_773 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_770 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_767 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_764 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_761 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_758 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_755 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_752 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_749 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_746 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_743 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_740 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_737 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_734 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_731 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_728 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_725 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_722 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_719 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_716 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_713 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_710 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_707 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_704 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_701 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_698 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_695 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_2139(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_2136(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2133(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2127(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2124(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2121(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2118(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2115(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2112(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2109(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2106(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2103(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2100(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2097(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2094(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(sum));
endmodule

module adder64__2_2284(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_2139 genblk1_48_F (.a(x[48]), .b(y[48]), .cin(), .sum(z[48]), .carry(
      carry[48]));
   FA__2_2136 genblk1_49_F (.a(x[49]), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(carry[49]));
   FA__2_2133 genblk1_50_F (.a(x[50]), .b(y[50]), .cin(carry[49]), .sum(z[50]), 
      .carry(carry[50]));
   FA__2_2130 genblk1_51_F (.a(x[51]), .b(y[51]), .cin(carry[50]), .sum(z[51]), 
      .carry(carry[51]));
   FA__2_2127 genblk1_52_F (.a(x[52]), .b(y[52]), .cin(carry[51]), .sum(z[52]), 
      .carry(carry[52]));
   FA__2_2124 genblk1_53_F (.a(x[53]), .b(y[53]), .cin(carry[52]), .sum(z[53]), 
      .carry(carry[53]));
   FA__2_2121 genblk1_54_F (.a(x[54]), .b(y[54]), .cin(carry[53]), .sum(z[54]), 
      .carry(carry[54]));
   FA__2_2118 genblk1_55_F (.a(x[55]), .b(y[55]), .cin(carry[54]), .sum(z[55]), 
      .carry(carry[55]));
   FA__2_2115 genblk1_56_F (.a(), .b(y[56]), .cin(carry[55]), .sum(z[56]), 
      .carry(carry[56]));
   FA__2_2112 genblk1_57_F (.a(), .b(y[57]), .cin(carry[56]), .sum(z[57]), 
      .carry(carry[57]));
   FA__2_2109 genblk1_58_F (.a(), .b(y[58]), .cin(carry[57]), .sum(z[58]), 
      .carry(carry[58]));
   FA__2_2106 genblk1_59_F (.a(), .b(y[59]), .cin(carry[58]), .sum(z[59]), 
      .carry(carry[59]));
   FA__2_2103 genblk1_60_F (.a(), .b(y[60]), .cin(carry[59]), .sum(z[60]), 
      .carry(carry[60]));
   FA__2_2100 genblk1_61_F (.a(), .b(y[61]), .cin(carry[60]), .sum(z[61]), 
      .carry(carry[61]));
   FA__2_2097 genblk1_62_F (.a(), .b(y[62]), .cin(carry[61]), .sum(z[62]), 
      .carry(carry[62]));
   FA__2_2094 genblk1_63_F (.a(), .b(y[63]), .cin(carry[62]), .sum(z[63]), 
      .carry());
endmodule

module FA__2_2356(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_2353(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2350(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2347(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2344(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2341(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2335(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2332(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2329(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2326(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2323(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2320(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2317(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2311(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2308(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2305(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2302(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2299(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2296(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2293(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2287(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(sum));
endmodule

module adder64__2_2477(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_2356 genblk1_40_F (.a(x[40]), .b(y[40]), .cin(), .sum(z[40]), .carry(
      carry[40]));
   FA__2_2353 genblk1_41_F (.a(x[41]), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__2_2350 genblk1_42_F (.a(x[42]), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__2_2347 genblk1_43_F (.a(x[43]), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__2_2344 genblk1_44_F (.a(x[44]), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__2_2341 genblk1_45_F (.a(x[45]), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__2_2338 genblk1_46_F (.a(x[46]), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__2_2335 genblk1_47_F (.a(x[47]), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__2_2332 genblk1_48_F (.a(x[48]), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(carry[48]));
   FA__2_2329 genblk1_49_F (.a(), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(carry[49]));
   FA__2_2326 genblk1_50_F (.a(), .b(y[50]), .cin(carry[49]), .sum(z[50]), 
      .carry(carry[50]));
   FA__2_2323 genblk1_51_F (.a(), .b(y[51]), .cin(carry[50]), .sum(z[51]), 
      .carry(carry[51]));
   FA__2_2320 genblk1_52_F (.a(), .b(y[52]), .cin(carry[51]), .sum(z[52]), 
      .carry(carry[52]));
   FA__2_2317 genblk1_53_F (.a(), .b(y[53]), .cin(carry[52]), .sum(z[53]), 
      .carry(carry[53]));
   FA__2_2314 genblk1_54_F (.a(), .b(y[54]), .cin(carry[53]), .sum(z[54]), 
      .carry(carry[54]));
   FA__2_2311 genblk1_55_F (.a(), .b(y[55]), .cin(carry[54]), .sum(z[55]), 
      .carry(carry[55]));
   FA__2_2308 genblk1_56_F (.a(), .b(y[56]), .cin(carry[55]), .sum(z[56]), 
      .carry(carry[56]));
   FA__2_2305 genblk1_57_F (.a(), .b(y[57]), .cin(carry[56]), .sum(z[57]), 
      .carry(carry[57]));
   FA__2_2302 genblk1_58_F (.a(), .b(y[58]), .cin(carry[57]), .sum(z[58]), 
      .carry(carry[58]));
   FA__2_2299 genblk1_59_F (.a(), .b(y[59]), .cin(carry[58]), .sum(z[59]), 
      .carry(carry[59]));
   FA__2_2296 genblk1_60_F (.a(), .b(y[60]), .cin(carry[59]), .sum(z[60]), 
      .carry(carry[60]));
   FA__2_2293 genblk1_61_F (.a(), .b(y[61]), .cin(carry[60]), .sum(z[61]), 
      .carry(carry[61]));
   FA__2_2290 genblk1_62_F (.a(), .b(y[62]), .cin(carry[61]), .sum(z[62]), 
      .carry(carry[62]));
   FA__2_2287 genblk1_63_F (.a(), .b(y[63]), .cin(carry[62]), .sum(z[63]), 
      .carry());
endmodule

module FA__2_2597(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_2594(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2591(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2588(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2585(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2582(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2579(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2576(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2573(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2567(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2564(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2561(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2558(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2555(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2552(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2549(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2546(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2543(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2540(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2537(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2534(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2531(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2528(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2525(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2519(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2516(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2513(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2510(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2507(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2504(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2501(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2495(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2492(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2489(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2486(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2483(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2480(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(sum));
endmodule

module adder64__2_2670(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_2597 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(), .sum(z[24]), .carry(
      carry[24]));
   FA__2_2594 genblk1_25_F (.a(x[25]), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__2_2591 genblk1_26_F (.a(x[26]), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__2_2588 genblk1_27_F (.a(x[27]), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__2_2585 genblk1_28_F (.a(x[28]), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__2_2582 genblk1_29_F (.a(x[29]), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__2_2579 genblk1_30_F (.a(x[30]), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__2_2576 genblk1_31_F (.a(x[31]), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__2_2573 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__2_2570 genblk1_33_F (.a(x[33]), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__2_2567 genblk1_34_F (.a(x[34]), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__2_2564 genblk1_35_F (.a(x[35]), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__2_2561 genblk1_36_F (.a(x[36]), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__2_2558 genblk1_37_F (.a(x[37]), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__2_2555 genblk1_38_F (.a(x[38]), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__2_2552 genblk1_39_F (.a(x[39]), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__2_2549 genblk1_40_F (.a(x[40]), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__2_2546 genblk1_41_F (.a(x[41]), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__2_2543 genblk1_42_F (.a(x[42]), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__2_2540 genblk1_43_F (.a(x[43]), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__2_2537 genblk1_44_F (.a(x[44]), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__2_2534 genblk1_45_F (.a(x[45]), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__2_2531 genblk1_46_F (.a(x[46]), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__2_2528 genblk1_47_F (.a(x[47]), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__2_2525 genblk1_48_F (.a(x[48]), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(carry[48]));
   FA__2_2522 genblk1_49_F (.a(x[49]), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(carry[49]));
   FA__2_2519 genblk1_50_F (.a(x[50]), .b(y[50]), .cin(carry[49]), .sum(z[50]), 
      .carry(carry[50]));
   FA__2_2516 genblk1_51_F (.a(x[51]), .b(y[51]), .cin(carry[50]), .sum(z[51]), 
      .carry(carry[51]));
   FA__2_2513 genblk1_52_F (.a(x[52]), .b(y[52]), .cin(carry[51]), .sum(z[52]), 
      .carry(carry[52]));
   FA__2_2510 genblk1_53_F (.a(x[53]), .b(y[53]), .cin(carry[52]), .sum(z[53]), 
      .carry(carry[53]));
   FA__2_2507 genblk1_54_F (.a(x[54]), .b(y[54]), .cin(carry[53]), .sum(z[54]), 
      .carry(carry[54]));
   FA__2_2504 genblk1_55_F (.a(x[55]), .b(y[55]), .cin(carry[54]), .sum(z[55]), 
      .carry(carry[55]));
   FA__2_2501 genblk1_56_F (.a(x[56]), .b(y[56]), .cin(carry[55]), .sum(z[56]), 
      .carry(carry[56]));
   FA__2_2498 genblk1_57_F (.a(x[57]), .b(y[57]), .cin(carry[56]), .sum(z[57]), 
      .carry(carry[57]));
   FA__2_2495 genblk1_58_F (.a(), .b(y[58]), .cin(carry[57]), .sum(z[58]), 
      .carry(carry[58]));
   FA__2_2492 genblk1_59_F (.a(), .b(y[59]), .cin(carry[58]), .sum(z[59]), 
      .carry(carry[59]));
   FA__2_2489 genblk1_60_F (.a(), .b(y[60]), .cin(carry[59]), .sum(z[60]), 
      .carry(carry[60]));
   FA__2_2486 genblk1_61_F (.a(), .b(y[61]), .cin(carry[60]), .sum(z[61]), 
      .carry(carry[61]));
   FA__2_2483 genblk1_62_F (.a(), .b(y[62]), .cin(carry[61]), .sum(z[62]), 
      .carry(carry[62]));
   FA__2_2480 genblk1_63_F (.a(), .b(y[63]), .cin(carry[62]), .sum(z[63]), 
      .carry());
endmodule

module FA__2_1135(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1132(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1129(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1126(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1123(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1120(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1117(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1111(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1108(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1105(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1102(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1099(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1096(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1093(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1090(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1087(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1084(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1081(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1078(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1075(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1072(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1069(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1066(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1063(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1060(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1057(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1054(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1051(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1048(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1045(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1042(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1039(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1036(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1033(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1030(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1027(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1024(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1021(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1015(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1012(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1009(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1006(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1003(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1000(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_997(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_991(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_988(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_985(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_982(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_979(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_976(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_973(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_970(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_967(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_964(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_961(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_958(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_955(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_952(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_949(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__2_1136(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_1135 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_1132 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_1129 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_1126 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_1123 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_1120 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_1117 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_1114 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_1111 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_1108 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_1105 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_1102 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_1099 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_1096 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_1093 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_1090 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_1087 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_1084 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_1081 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_1078 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_1075 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_1072 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_1069 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_1066 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_1063 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_1060 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_1057 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_1054 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_1051 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_1048 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_1045 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_1042 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_1039 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_1036 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_1033 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_1030 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_1027 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_1024 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_1021 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_1018 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_1015 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_1012 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_1009 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_1006 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_1003 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_1000 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_997 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_994 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_991 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_988 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_985 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_982 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_979 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_976 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_973 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_970 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_967 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_964 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_961 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_958 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_955 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_952 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_949 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_2766(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_2763(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2760(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2757(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2751(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2748(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2745(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2742(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2739(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2736(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2733(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2727(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2724(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2721(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2718(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2715(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2712(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2709(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2703(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2700(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2697(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2694(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__2_2863(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_2766 genblk1_32_F (.a(x[32]), .b(y[32]), .cin(), .sum(z[32]), .carry(
      carry[32]));
   FA__2_2763 genblk1_33_F (.a(x[33]), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__2_2760 genblk1_34_F (.a(x[34]), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__2_2757 genblk1_35_F (.a(x[35]), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__2_2754 genblk1_36_F (.a(x[36]), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__2_2751 genblk1_37_F (.a(x[37]), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__2_2748 genblk1_38_F (.a(x[38]), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__2_2745 genblk1_39_F (.a(x[39]), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(carry[39]));
   FA__2_2742 genblk1_40_F (.a(x[40]), .b(y[40]), .cin(carry[39]), .sum(z[40]), 
      .carry(carry[40]));
   FA__2_2739 genblk1_41_F (.a(), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__2_2736 genblk1_42_F (.a(), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__2_2733 genblk1_43_F (.a(), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__2_2730 genblk1_44_F (.a(), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__2_2727 genblk1_45_F (.a(), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__2_2724 genblk1_46_F (.a(), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__2_2721 genblk1_47_F (.a(), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__2_2718 genblk1_48_F (.a(), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(carry[48]));
   FA__2_2715 genblk1_49_F (.a(), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(carry[49]));
   FA__2_2712 genblk1_50_F (.a(), .b(y[50]), .cin(carry[49]), .sum(z[50]), 
      .carry(carry[50]));
   FA__2_2709 genblk1_51_F (.a(), .b(y[51]), .cin(carry[50]), .sum(z[51]), 
      .carry(carry[51]));
   FA__2_2706 genblk1_52_F (.a(), .b(y[52]), .cin(carry[51]), .sum(z[52]), 
      .carry(carry[52]));
   FA__2_2703 genblk1_53_F (.a(), .b(y[53]), .cin(carry[52]), .sum(z[53]), 
      .carry(carry[53]));
   FA__2_2700 genblk1_54_F (.a(), .b(y[54]), .cin(carry[53]), .sum(z[54]), 
      .carry(carry[54]));
   FA__2_2697 genblk1_55_F (.a(), .b(y[55]), .cin(carry[54]), .sum(z[55]), 
      .carry(carry[55]));
   FA__2_2694 genblk1_56_F (.a(), .b(y[56]), .cin(carry[55]), .sum(z[56]), 
      .carry(z[57]));
endmodule

module FA__2_2935(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_2932(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2929(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2926(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2923(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2920(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2917(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2914(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_2911(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2908(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2905(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2902(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2899(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2896(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2893(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_2890(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64__2_3056(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_2935 genblk1_40_F (.a(x[40]), .b(y[40]), .cin(), .sum(z[40]), .carry(
      carry[40]));
   FA__2_2932 genblk1_41_F (.a(x[41]), .b(y[41]), .cin(carry[40]), .sum(z[41]), 
      .carry(carry[41]));
   FA__2_2929 genblk1_42_F (.a(x[42]), .b(y[42]), .cin(carry[41]), .sum(z[42]), 
      .carry(carry[42]));
   FA__2_2926 genblk1_43_F (.a(x[43]), .b(y[43]), .cin(carry[42]), .sum(z[43]), 
      .carry(carry[43]));
   FA__2_2923 genblk1_44_F (.a(x[44]), .b(y[44]), .cin(carry[43]), .sum(z[44]), 
      .carry(carry[44]));
   FA__2_2920 genblk1_45_F (.a(x[45]), .b(y[45]), .cin(carry[44]), .sum(z[45]), 
      .carry(carry[45]));
   FA__2_2917 genblk1_46_F (.a(x[46]), .b(y[46]), .cin(carry[45]), .sum(z[46]), 
      .carry(carry[46]));
   FA__2_2914 genblk1_47_F (.a(x[47]), .b(y[47]), .cin(carry[46]), .sum(z[47]), 
      .carry(carry[47]));
   FA__2_2911 genblk1_48_F (.a(), .b(y[48]), .cin(carry[47]), .sum(z[48]), 
      .carry(carry[48]));
   FA__2_2908 genblk1_49_F (.a(), .b(y[49]), .cin(carry[48]), .sum(z[49]), 
      .carry(carry[49]));
   FA__2_2905 genblk1_50_F (.a(), .b(y[50]), .cin(carry[49]), .sum(z[50]), 
      .carry(carry[50]));
   FA__2_2902 genblk1_51_F (.a(), .b(y[51]), .cin(carry[50]), .sum(z[51]), 
      .carry(carry[51]));
   FA__2_2899 genblk1_52_F (.a(), .b(y[52]), .cin(carry[51]), .sum(z[52]), 
      .carry(carry[52]));
   FA__2_2896 genblk1_53_F (.a(), .b(y[53]), .cin(carry[52]), .sum(z[53]), 
      .carry(carry[53]));
   FA__2_2893 genblk1_54_F (.a(), .b(y[54]), .cin(carry[53]), .sum(z[54]), 
      .carry(carry[54]));
   FA__2_2890 genblk1_55_F (.a(), .b(y[55]), .cin(carry[54]), .sum(z[55]), 
      .carry(z[56]));
endmodule

module FA__2_1389(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1383(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1380(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1377(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1374(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1371(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1368(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1365(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1359(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1356(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1353(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1350(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1347(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1344(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1341(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1335(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1332(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1329(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1326(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1323(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1320(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1317(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1311(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1308(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1305(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1302(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1299(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1296(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1293(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1287(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1284(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1281(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1278(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1275(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1272(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1269(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1263(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1260(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1257(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1254(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1251(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1248(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1245(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1242(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1239(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1236(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1233(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1230(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1227(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1224(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1221(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1215(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1212(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1209(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1206(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1203(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__2_1390(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_1389 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_1386 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_1383 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_1380 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_1377 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_1374 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_1371 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_1368 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_1365 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_1362 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_1359 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_1356 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_1353 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_1350 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_1347 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_1344 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_1341 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_1338 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_1335 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_1332 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_1329 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_1326 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_1323 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_1320 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_1317 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_1314 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_1311 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_1308 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_1305 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_1302 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_1299 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_1296 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_1293 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_1290 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_1287 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_1284 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_1281 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_1278 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_1275 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_1272 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_1269 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_1266 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_1263 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_1260 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_1257 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_1254 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_1251 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_1248 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_1245 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_1242 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_1239 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_1236 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_1233 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_1230 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_1227 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_1224 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_1221 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_1218 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_1215 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_1212 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_1209 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_1206 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_1203 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_212(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(carry));
endmodule

module FA__2_215(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_221(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_224(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_227(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_230(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_233(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_236(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_239(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_245(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_248(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_251(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_254(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module FA__2_257(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(cin), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(carry));
endmodule

module adder64(x, y, z, C);
   input [63:0]x;
   input [63:0]y;
   output [63:0]z;
   output C;

   wire [64:0]carry;

   FA__2_212 genblk1_24_F (.a(x[24]), .b(y[24]), .cin(), .sum(z[24]), .carry(
      carry[24]));
   FA__2_215 genblk1_25_F (.a(x[25]), .b(y[25]), .cin(carry[24]), .sum(z[25]), 
      .carry(carry[25]));
   FA__2_218 genblk1_26_F (.a(x[26]), .b(y[26]), .cin(carry[25]), .sum(z[26]), 
      .carry(carry[26]));
   FA__2_221 genblk1_27_F (.a(x[27]), .b(y[27]), .cin(carry[26]), .sum(z[27]), 
      .carry(carry[27]));
   FA__2_224 genblk1_28_F (.a(x[28]), .b(y[28]), .cin(carry[27]), .sum(z[28]), 
      .carry(carry[28]));
   FA__2_227 genblk1_29_F (.a(x[29]), .b(y[29]), .cin(carry[28]), .sum(z[29]), 
      .carry(carry[29]));
   FA__2_230 genblk1_30_F (.a(x[30]), .b(y[30]), .cin(carry[29]), .sum(z[30]), 
      .carry(carry[30]));
   FA__2_233 genblk1_31_F (.a(x[31]), .b(y[31]), .cin(carry[30]), .sum(z[31]), 
      .carry(carry[31]));
   FA__2_236 genblk1_32_F (.a(), .b(y[32]), .cin(carry[31]), .sum(z[32]), 
      .carry(carry[32]));
   FA__2_239 genblk1_33_F (.a(), .b(y[33]), .cin(carry[32]), .sum(z[33]), 
      .carry(carry[33]));
   FA__2_242 genblk1_34_F (.a(), .b(y[34]), .cin(carry[33]), .sum(z[34]), 
      .carry(carry[34]));
   FA__2_245 genblk1_35_F (.a(), .b(y[35]), .cin(carry[34]), .sum(z[35]), 
      .carry(carry[35]));
   FA__2_248 genblk1_36_F (.a(), .b(y[36]), .cin(carry[35]), .sum(z[36]), 
      .carry(carry[36]));
   FA__2_251 genblk1_37_F (.a(), .b(y[37]), .cin(carry[36]), .sum(z[37]), 
      .carry(carry[37]));
   FA__2_254 genblk1_38_F (.a(), .b(y[38]), .cin(carry[37]), .sum(z[38]), 
      .carry(carry[38]));
   FA__2_257 genblk1_39_F (.a(), .b(y[39]), .cin(carry[38]), .sum(z[39]), 
      .carry(z[40]));
endmodule

module FA__2_1643(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1640(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1637(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1634(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1631(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1628(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1625(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1622(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1619(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1616(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1613(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1610(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1607(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1604(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1601(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1598(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1595(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1592(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1589(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1586(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1583(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1580(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1577(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1574(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1571(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1568(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1565(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1559(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1556(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1553(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1550(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1547(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1544(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1541(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1538(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1535(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1532(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1529(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1526(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1523(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1520(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1517(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1511(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1508(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1505(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1502(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1499(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1496(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1493(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1490(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1487(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1484(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1481(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1478(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1475(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1472(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1469(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1463(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1460(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1457(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__2_1644(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_1643 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_1640 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_1637 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_1634 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_1631 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_1628 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_1625 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_1622 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_1619 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_1616 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_1613 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_1610 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_1607 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_1604 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_1601 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_1598 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_1595 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_1592 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_1589 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_1586 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_1583 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_1580 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_1577 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_1574 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_1571 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_1568 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_1565 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_1562 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_1559 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_1556 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_1553 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_1550 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_1547 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_1544 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_1541 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_1538 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_1535 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_1532 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_1529 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_1526 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_1523 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_1520 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_1517 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_1514 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_1511 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_1508 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_1505 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_1502 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_1499 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_1496 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_1493 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_1490 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_1487 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_1484 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_1481 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_1478 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_1475 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_1472 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_1469 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_1466 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_1463 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_1460 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_1457 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_1897(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1894(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1891(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1888(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1885(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1882(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1879(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1876(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1873(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1870(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1867(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1864(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1861(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1858(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1855(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1852(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_1849(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1846(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1843(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1840(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1837(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1831(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1828(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1825(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1822(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1819(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1816(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1813(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1807(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1804(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1801(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1798(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1795(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1792(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1789(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1783(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1780(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1777(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1774(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1771(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1768(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1765(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1759(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1756(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1753(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1750(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1747(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1744(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1741(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1735(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1732(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1729(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1726(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1723(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1720(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_1717(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_1714(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_1711(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8__2_1898(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_1897 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_1894 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_1891 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_1888 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_1885 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_1882 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_1879 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_1876 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_1873 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_1870 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_1867 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_1864 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_1861 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_1858 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_1855 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_1852 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_1849 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_1846 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_1843 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_1840 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_1837 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_1834 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_1831 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_1828 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_1825 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_1822 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_1819 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_1816 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_1813 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_1810 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_1807 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_1804 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_1801 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_1798 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_1795 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_1792 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_1789 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_1786 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_1783 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_1780 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_1777 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_1774 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_1771 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_1768 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_1765 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_1762 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_1759 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_1756 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_1753 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_1750 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_1747 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_1744 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_1741 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_1738 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_1735 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_1732 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_1729 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_1726 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_1723 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_1720 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_1717 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_1714 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_1711 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module FA__2_2(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_5(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_8(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_11(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_14(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_329(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_17(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_20(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_23(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_26(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_332(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_335(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_338(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_341(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_344(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_347(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module HA__2_350(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_29(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_32(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_35(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_353(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_38(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_356(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_41(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_44(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_47(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_50(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_53(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_56(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_59(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_62(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_359(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_65(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_68(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_71(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_74(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_77(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_80(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_83(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_86(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_89(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_92(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_95(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_98(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_101(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_104(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_107(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_110(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_113(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_362(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_116(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_365(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_119(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_122(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_125(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_368(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_128(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_131(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_371(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_134(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module FA__2_137(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(carry));
   OAI21_X1 i_0_1 (.A(b), .B1(cin), .B2(a), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(b), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(a), .ZN(n_0_2));
endmodule

module HA__2_374(a, b, s, c);
   input a;
   input b;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(s));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(c));
endmodule

module FA__2_140(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(a), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(b), .ZN(sum));
endmodule

module WTM8(A, B, Result);
   input [7:0]A;
   input [7:0]B;
   output [15:0]Result;

   wire C;
   wire S;
   wire P;

   FA__2_2 F3 (.a(n_155), .b(n_147), .cin(n_139), .sum(S), .carry(C));
   FA__2_5 F2 (.a(n_161), .b(n_154), .cin(n_146), .sum(n_1), .carry(n_0));
   FA__2_8 F7 (.a(n_131), .b(n_123), .cin(n_116), .sum(n_3), .carry(n_2));
   FA__2_11 F14 (.a(S), .b(n_0), .cin(n_3), .sum(n_5), .carry(n_4));
   FA__2_14 F1 (.a(n_160), .b(n_153), .cin(n_145), .sum(n_7), .carry(n_6));
   HA__2_329 H2 (.a(n_138), .b(n_130), .s(n_9), .c(n_8));
   FA__2_17 F13 (.a(n_1), .b(n_6), .cin(n_9), .sum(n_11), .carry(n_10));
   FA__2_20 F25 (.a(n_5), .b(n_10), .cin(n_8), .sum(n_13), .carry(n_12));
   FA__2_23 F0 (.a(n_159), .b(n_152), .cin(n_144), .sum(n_15), .carry(n_14));
   FA__2_26 F12 (.a(n_7), .b(n_14), .cin(n_137), .sum(n_17), .carry(n_16));
   HA__2_332 H8 (.a(n_11), .b(n_16), .s(n_19), .c(n_18));
   HA__2_335 H12 (.a(n_13), .b(n_18), .s(n_21), .c(n_20));
   HA__2_338 H0 (.a(n_158), .b(n_151), .s(Result[1]), .c(n_22));
   HA__2_341 H4 (.a(n_15), .b(n_22), .s(Result[2]), .c(n_23));
   HA__2_344 H7 (.a(n_17), .b(n_23), .s(Result[3]), .c(n_24));
   HA__2_347 H11 (.a(n_19), .b(n_24), .s(Result[4]), .c(n_25));
   HA__2_350 H15 (.a(n_21), .b(n_25), .s(Result[5]), .c(n_26));
   FA__2_29 F4 (.a(n_156), .b(n_148), .cin(n_140), .sum(n_28), .carry(n_27));
   FA__2_32 F8 (.a(n_132), .b(n_124), .cin(n_117), .sum(n_30), .carry(n_29));
   FA__2_35 F15 (.a(n_28), .b(C), .cin(n_30), .sum(n_32), .carry(n_31));
   HA__2_353 H6 (.a(n_162), .b(n_2), .s(n_34), .c(n_33));
   FA__2_38 F26 (.a(n_32), .b(n_4), .cin(n_34), .sum(n_36), .carry(n_35));
   HA__2_356 H13 (.a(n_36), .b(n_12), .s(n_38), .c(n_37));
   FA__2_41 F38 (.a(n_38), .b(n_20), .cin(n_26), .sum(Result[6]), .carry(n_39));
   FA__2_44 F5 (.a(n_157), .b(n_149), .cin(n_141), .sum(n_41), .carry(n_40));
   FA__2_47 F9 (.a(n_133), .b(n_125), .cin(n_118), .sum(n_43), .carry(n_42));
   FA__2_50 F16 (.a(n_41), .b(n_27), .cin(n_43), .sum(n_45), .carry(n_44));
   FA__2_53 F22 (.a(n_29), .b(n_163), .cin(n_108), .sum(n_47), .carry(n_46));
   FA__2_56 F27 (.a(n_45), .b(n_31), .cin(n_47), .sum(n_49), .carry(n_48));
   FA__2_59 F31 (.a(n_49), .b(n_35), .cin(n_33), .sum(n_51), .carry(n_50));
   FA__2_62 F39 (.a(n_51), .b(n_37), .cin(n_39), .sum(Result[7]), .carry(n_52));
   HA__2_359 H1 (.a(n_150), .b(n_142), .s(n_54), .c(n_53));
   FA__2_65 F10 (.a(n_134), .b(n_126), .cin(n_120), .sum(n_56), .carry(n_55));
   FA__2_68 F17 (.a(n_54), .b(n_40), .cin(n_56), .sum(n_58), .carry(n_57));
   FA__2_71 F23 (.a(n_42), .b(n_164), .cin(n_109), .sum(n_60), .carry(n_59));
   FA__2_74 F28 (.a(n_58), .b(n_44), .cin(n_60), .sum(n_62), .carry(n_61));
   FA__2_77 F32 (.a(n_62), .b(n_48), .cin(n_46), .sum(n_64), .carry(n_63));
   FA__2_80 F40 (.a(n_64), .b(n_50), .cin(n_52), .sum(Result[8]), .carry(n_65));
   FA__2_83 F6 (.a(n_143), .b(n_135), .cin(n_127), .sum(n_67), .carry(n_66));
   FA__2_86 F18 (.a(n_67), .b(n_53), .cin(n_55), .sum(n_69), .carry(n_68));
   FA__2_89 F24 (.a(n_119), .b(n_165), .cin(n_110), .sum(n_71), .carry(n_70));
   FA__2_92 F29 (.a(n_69), .b(n_57), .cin(n_71), .sum(n_73), .carry(n_72));
   FA__2_95 F33 (.a(n_73), .b(n_61), .cin(n_59), .sum(n_75), .carry(n_74));
   FA__2_98 F41 (.a(n_75), .b(n_63), .cin(n_65), .sum(Result[9]), .carry(n_76));
   FA__2_101 F11 (.a(n_136), .b(n_128), .cin(n_121), .sum(n_78), .carry(n_77));
   FA__2_104 F19 (.a(n_66), .b(n_166), .cin(n_111), .sum(n_80), .carry(n_79));
   FA__2_107 F30 (.a(n_78), .b(n_68), .cin(n_80), .sum(n_82), .carry(n_81));
   FA__2_110 F34 (.a(n_82), .b(n_72), .cin(n_70), .sum(n_84), .carry(n_83));
   FA__2_113 F42 (.a(n_84), .b(n_74), .cin(n_76), .sum(Result[10]), .carry(n_85));
   HA__2_362 H3 (.a(n_129), .b(P), .s(n_87), .c(n_86));
   FA__2_116 F20 (.a(n_77), .b(n_167), .cin(n_112), .sum(n_89), .carry(n_88));
   HA__2_365 H9 (.a(n_87), .b(n_89), .s(n_91), .c(n_90));
   FA__2_119 F35 (.a(n_91), .b(n_81), .cin(n_79), .sum(n_93), .carry(n_92));
   FA__2_122 F43 (.a(n_93), .b(n_83), .cin(n_85), .sum(Result[11]), .carry(n_94));
   FA__2_125 F21 (.a(n_122), .b(n_168), .cin(n_113), .sum(n_96), .carry(n_95));
   HA__2_368 H10 (.a(n_86), .b(n_96), .s(n_98), .c(n_97));
   FA__2_128 F36 (.a(n_98), .b(n_88), .cin(n_90), .sum(n_100), .carry(n_99));
   FA__2_131 F44 (.a(n_100), .b(n_92), .cin(n_94), .sum(Result[12]), .carry(
      n_101));
   HA__2_371 H5 (.a(n_169), .b(n_114), .s(n_103), .c(n_102));
   FA__2_134 F37 (.a(n_97), .b(n_103), .cin(n_95), .sum(n_105), .carry(n_104));
   FA__2_137 F45 (.a(n_105), .b(n_99), .cin(n_101), .sum(Result[13]), .carry(
      n_106));
   HA__2_374 H14 (.a(n_115), .b(n_102), .s(n_107), .c(Result[15]));
   FA__2_140 F46 (.a(n_107), .b(n_104), .cin(n_106), .sum(Result[14]), .carry());
   AND2_X1 i_0_0 (.A1(A[0]), .A2(B[0]), .ZN(Result[0]));
   AND2_X1 i_0_1 (.A1(A[0]), .A2(B[7]), .ZN(n_108));
   AND2_X1 i_0_2 (.A1(A[1]), .A2(B[7]), .ZN(n_109));
   AND2_X1 i_0_3 (.A1(A[2]), .A2(B[7]), .ZN(n_110));
   AND2_X1 i_0_4 (.A1(A[3]), .A2(B[7]), .ZN(n_111));
   AND2_X1 i_0_5 (.A1(A[4]), .A2(B[7]), .ZN(n_112));
   AND2_X1 i_0_6 (.A1(A[5]), .A2(B[7]), .ZN(n_113));
   AND2_X1 i_0_7 (.A1(A[6]), .A2(B[7]), .ZN(n_114));
   AND2_X1 i_0_8 (.A1(A[7]), .A2(B[7]), .ZN(n_115));
   AND2_X1 i_0_9 (.A1(A[0]), .A2(B[5]), .ZN(n_116));
   AND2_X1 i_0_10 (.A1(A[1]), .A2(B[5]), .ZN(n_117));
   AND2_X1 i_0_11 (.A1(A[2]), .A2(B[5]), .ZN(n_118));
   AND2_X1 i_0_12 (.A1(A[4]), .A2(B[5]), .ZN(n_119));
   AND2_X1 i_0_13 (.A1(A[3]), .A2(B[5]), .ZN(n_120));
   AND2_X1 i_0_14 (.A1(A[5]), .A2(B[5]), .ZN(n_121));
   AND2_X1 i_0_15 (.A1(A[7]), .A2(B[5]), .ZN(n_122));
   AND2_X1 i_0_16 (.A1(A[6]), .A2(B[5]), .ZN(P));
   AND2_X1 i_0_17 (.A1(A[1]), .A2(B[4]), .ZN(n_123));
   AND2_X1 i_0_18 (.A1(A[2]), .A2(B[4]), .ZN(n_124));
   AND2_X1 i_0_19 (.A1(A[3]), .A2(B[4]), .ZN(n_125));
   AND2_X1 i_0_20 (.A1(A[4]), .A2(B[4]), .ZN(n_126));
   AND2_X1 i_0_21 (.A1(A[5]), .A2(B[4]), .ZN(n_127));
   AND2_X1 i_0_22 (.A1(A[6]), .A2(B[4]), .ZN(n_128));
   AND2_X1 i_0_23 (.A1(A[7]), .A2(B[4]), .ZN(n_129));
   AND2_X1 i_0_24 (.A1(A[0]), .A2(B[4]), .ZN(n_130));
   AND2_X1 i_0_25 (.A1(A[2]), .A2(B[3]), .ZN(n_131));
   AND2_X1 i_0_26 (.A1(A[3]), .A2(B[3]), .ZN(n_132));
   AND2_X1 i_0_27 (.A1(A[4]), .A2(B[3]), .ZN(n_133));
   AND2_X1 i_0_28 (.A1(A[5]), .A2(B[3]), .ZN(n_134));
   AND2_X1 i_0_29 (.A1(A[6]), .A2(B[3]), .ZN(n_135));
   AND2_X1 i_0_30 (.A1(A[7]), .A2(B[3]), .ZN(n_136));
   AND2_X1 i_0_31 (.A1(A[0]), .A2(B[3]), .ZN(n_137));
   AND2_X1 i_0_32 (.A1(A[1]), .A2(B[3]), .ZN(n_138));
   AND2_X1 i_0_33 (.A1(A[3]), .A2(B[2]), .ZN(n_139));
   AND2_X1 i_0_34 (.A1(A[4]), .A2(B[2]), .ZN(n_140));
   AND2_X1 i_0_35 (.A1(A[5]), .A2(B[2]), .ZN(n_141));
   AND2_X1 i_0_36 (.A1(A[6]), .A2(B[2]), .ZN(n_142));
   AND2_X1 i_0_37 (.A1(A[7]), .A2(B[2]), .ZN(n_143));
   AND2_X1 i_0_38 (.A1(A[0]), .A2(B[2]), .ZN(n_144));
   AND2_X1 i_0_39 (.A1(A[1]), .A2(B[2]), .ZN(n_145));
   AND2_X1 i_0_40 (.A1(A[2]), .A2(B[2]), .ZN(n_146));
   AND2_X1 i_0_41 (.A1(A[4]), .A2(B[1]), .ZN(n_147));
   AND2_X1 i_0_42 (.A1(A[5]), .A2(B[1]), .ZN(n_148));
   AND2_X1 i_0_43 (.A1(A[6]), .A2(B[1]), .ZN(n_149));
   AND2_X1 i_0_44 (.A1(A[7]), .A2(B[1]), .ZN(n_150));
   AND2_X1 i_0_45 (.A1(A[0]), .A2(B[1]), .ZN(n_151));
   AND2_X1 i_0_46 (.A1(A[1]), .A2(B[1]), .ZN(n_152));
   AND2_X1 i_0_47 (.A1(A[2]), .A2(B[1]), .ZN(n_153));
   AND2_X1 i_0_48 (.A1(A[3]), .A2(B[1]), .ZN(n_154));
   AND2_X1 i_0_49 (.A1(A[5]), .A2(B[0]), .ZN(n_155));
   AND2_X1 i_0_50 (.A1(A[6]), .A2(B[0]), .ZN(n_156));
   AND2_X1 i_0_51 (.A1(A[7]), .A2(B[0]), .ZN(n_157));
   AND2_X1 i_0_52 (.A1(A[1]), .A2(B[0]), .ZN(n_158));
   AND2_X1 i_0_53 (.A1(A[2]), .A2(B[0]), .ZN(n_159));
   AND2_X1 i_0_54 (.A1(A[3]), .A2(B[0]), .ZN(n_160));
   AND2_X1 i_0_55 (.A1(A[4]), .A2(B[0]), .ZN(n_161));
   AND2_X1 i_0_56 (.A1(A[0]), .A2(B[6]), .ZN(n_162));
   AND2_X1 i_0_57 (.A1(A[1]), .A2(B[6]), .ZN(n_163));
   AND2_X1 i_0_58 (.A1(A[2]), .A2(B[6]), .ZN(n_164));
   AND2_X1 i_0_59 (.A1(A[3]), .A2(B[6]), .ZN(n_165));
   AND2_X1 i_0_60 (.A1(A[4]), .A2(B[6]), .ZN(n_166));
   AND2_X1 i_0_61 (.A1(A[5]), .A2(B[6]), .ZN(n_167));
   AND2_X1 i_0_62 (.A1(A[6]), .A2(B[6]), .ZN(n_168));
   AND2_X1 i_0_63 (.A1(A[7]), .A2(B[6]), .ZN(n_169));
endmodule

module WTM32(A, B, Result);
   input [31:0]A;
   input [31:0]B;
   output [63:0]Result;

   wire [15:0]\P[0] ;
   wire [63:0]\couple[0] ;
   wire [15:0]\P[2] ;
   wire [15:0]\P[3] ;
   wire [63:0]\couple[1] ;
   wire [63:0]\Quadruple[0] ;
   wire [15:0]\P[4] ;
   wire [15:0]\P[5] ;
   wire [63:0]\couple[2] ;
   wire [15:0]\P[6] ;
   wire [15:0]\P[7] ;
   wire [63:0]\couple[3] ;
   wire [63:0]\Quadruple[1] ;
   wire [63:0]\Eight[0] ;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire [15:0]\P[10] ;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_62;
   wire [63:0]out;
   wire [15:0]\P[14] ;
   wire [31:0]b;
   wire [31:0]a;
   wire n_0_0_0;
   wire [63:0]\couple[6] ;
   wire [15:0]\P[13] ;
   wire [15:0]\P[15] ;
   wire [63:0]\couple[7] ;
   wire [63:0]\Quadruple[3] ;
   wire [63:0]\Eight[1] ;
   wire [15:0]\P[12] ;
   wire [63:0]\Quadruple[2] ;
   wire [63:0]\couple[5] ;
   wire [15:0]\P[11] ;
   wire [63:0]\couple[4] ;
   wire [15:0]\P[9] ;
   wire [15:0]\P[8] ;
   wire [15:0]\P[1] ;

   WTM8__1_628 M0 (.A({a[7], a[6], a[5], a[4], a[3], a[2], a[1], A[0]}), 
      .B({b[7], b[6], b[5], b[4], b[3], b[2], b[1], B[0]}), .Result({\P[0] [15], 
      \P[0] [14], \P[0] [13], \P[0] [12], \P[0] [11], \P[0] [10], \P[0] [9], 
      \P[0] [8], \P[0] [7], \P[0] [6], \P[0] [5], \P[0] [4], \P[0] [3], 
      \P[0] [2], \P[0] [1], Result[0]}));
   adder64__1_2599 A0 (.x({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, 
      uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, 
      uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, \P[0] [15], 
      \P[0] [14], \P[0] [13], \P[0] [12], \P[0] [11], \P[0] [10], \P[0] [9], 
      \P[0] [8], uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55}), 
      .y({uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, 
      uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, 
      uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, 
      uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, 
      \P[1] [15], \P[1] [14], \P[1] [13], \P[1] [12], \P[1] [11], \P[1] [10], 
      \P[1] [9], \P[1] [8], \P[1] [7], \P[1] [6], \P[1] [5], \P[1] [4], 
      \P[1] [3], \P[1] [2], \P[1] [1], \P[1] [0], uc_96, uc_97, uc_98, uc_99, 
      uc_100, uc_101, uc_102, uc_103}), .z({uc_104, uc_105, uc_106, uc_107, 
      uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, 
      uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, 
      uc_126, uc_127, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, 
      uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, 
      \couple[0] [24], \couple[0] [23], \couple[0] [22], \couple[0] [21], 
      \couple[0] [20], \couple[0] [19], \couple[0] [18], \couple[0] [17], 
      \couple[0] [16], \couple[0] [15], \couple[0] [14], \couple[0] [13], 
      \couple[0] [12], \couple[0] [11], \couple[0] [10], \couple[0] [9], 
      \couple[0] [8], uc_143, uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, 
      uc_150}), .C());
   WTM8__1_882 M2 (.A({a[7], a[6], a[5], a[4], a[3], a[2], a[1], A[0]}), 
      .B({b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16]}), .Result(
      \P[2] ));
   WTM8__1_1136 M3 (.A({a[7], a[6], a[5], a[4], a[3], a[2], a[1], A[0]}), 
      .B({b[31], b[30], b[29], b[28], b[27], b[26], b[25], b[24]}), .Result(
      \P[3] ));
   adder64__1_2792 A1 (.x({uc_151, uc_152, uc_153, uc_154, uc_155, uc_156, 
      uc_157, uc_158, uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, 
      uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, 
      uc_175, uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, \P[2] [15], 
      \P[2] [14], \P[2] [13], \P[2] [12], \P[2] [11], \P[2] [10], \P[2] [9], 
      \P[2] [8], uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, uc_189, uc_190, 
      uc_191, uc_192, uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, 
      uc_200, uc_201, uc_202, uc_203, uc_204, uc_205, uc_206}), .y({uc_207, 
      uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, uc_216, 
      uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, uc_225, 
      uc_226, uc_227, uc_228, uc_229, uc_230, \P[3] [15], \P[3] [14], \P[3] [13], 
      \P[3] [12], \P[3] [11], \P[3] [10], \P[3] [9], \P[3] [8], \P[3] [7], 
      \P[3] [6], \P[3] [5], \P[3] [4], \P[3] [3], \P[3] [2], \P[3] [1], 
      \P[3] [0], uc_231, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, 
      uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, 
      uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254}), .z({uc_255, 
      uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, uc_262, uc_263, uc_264, 
      uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, 
      uc_274, uc_275, uc_276, uc_277, \couple[1] [40], \couple[1] [39], 
      \couple[1] [38], \couple[1] [37], \couple[1] [36], \couple[1] [35], 
      \couple[1] [34], \couple[1] [33], \couple[1] [32], \couple[1] [31], 
      \couple[1] [30], \couple[1] [29], \couple[1] [28], \couple[1] [27], 
      \couple[1] [26], \couple[1] [25], \couple[1] [24], uc_278, uc_279, uc_280, 
      uc_281, uc_282, uc_283, uc_284, uc_285, uc_286, uc_287, uc_288, uc_289, 
      uc_290, uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297, uc_298, 
      uc_299, uc_300, uc_301}), .C());
   adder64__1_2985 A8 (.x({uc_302, uc_303, uc_304, uc_305, uc_306, uc_307, 
      uc_308, uc_309, uc_310, uc_311, uc_312, uc_313, uc_314, uc_315, uc_316, 
      uc_317, uc_318, uc_319, uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, 
      uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, uc_334, 
      uc_335, uc_336, uc_337, uc_338, uc_339, uc_340, \couple[0] [24], 
      \couple[0] [23], \couple[0] [22], \couple[0] [21], \couple[0] [20], 
      \couple[0] [19], \couple[0] [18], \couple[0] [17], \couple[0] [16], uc_341, 
      uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, uc_348, uc_349, uc_350, 
      uc_351, uc_352, uc_353, uc_354, uc_355, uc_356}), .y({uc_357, uc_358, 
      uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, uc_366, uc_367, 
      uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, uc_376, 
      uc_377, uc_378, uc_379, \couple[1] [40], \couple[1] [39], \couple[1] [38], 
      \couple[1] [37], \couple[1] [36], \couple[1] [35], \couple[1] [34], 
      \couple[1] [33], \couple[1] [32], \couple[1] [31], \couple[1] [30], 
      \couple[1] [29], \couple[1] [28], \couple[1] [27], \couple[1] [26], 
      \couple[1] [25], \couple[1] [24], \P[2] [7], \P[2] [6], \P[2] [5], 
      \P[2] [4], \P[2] [3], \P[2] [2], \P[2] [1], \P[2] [0], uc_380, uc_381, 
      uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, 
      uc_391, uc_392, uc_393, uc_394, uc_395}), .z({uc_396, uc_397, uc_398, 
      uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, 
      uc_408, uc_409, uc_410, uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, 
      uc_417, \Quadruple[0] [41], \Quadruple[0] [40], \Quadruple[0] [39], 
      \Quadruple[0] [38], \Quadruple[0] [37], \Quadruple[0] [36], 
      \Quadruple[0] [35], \Quadruple[0] [34], \Quadruple[0] [33], 
      \Quadruple[0] [32], \Quadruple[0] [31], \Quadruple[0] [30], 
      \Quadruple[0] [29], \Quadruple[0] [28], \Quadruple[0] [27], 
      \Quadruple[0] [26], \Quadruple[0] [25], \Quadruple[0] [24], 
      \Quadruple[0] [23], \Quadruple[0] [22], \Quadruple[0] [21], 
      \Quadruple[0] [20], \Quadruple[0] [19], \Quadruple[0] [18], 
      \Quadruple[0] [17], \Quadruple[0] [16], uc_418, uc_419, uc_420, uc_421, 
      uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, uc_430, 
      uc_431, uc_432, uc_433}), .C());
   WTM8__1_1390 M4 (.A({a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8]}), 
      .B({b[7], b[6], b[5], b[4], b[3], b[2], b[1], B[0]}), .Result(\P[4] ));
   WTM8__1_1644 M5 (.A({a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8]}), 
      .B({b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8]}), .Result(\P[5] ));
   adder64__1_3178 A2 (.x({uc_434, uc_435, uc_436, uc_437, uc_438, uc_439, 
      uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, 
      uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, 
      uc_458, uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, uc_465, uc_466, 
      uc_467, uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, \P[4] [15], 
      \P[4] [14], \P[4] [13], \P[4] [12], \P[4] [11], \P[4] [10], \P[4] [9], 
      \P[4] [8], uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, 
      uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489}), .y({
      uc_490, uc_491, uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, 
      uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, 
      uc_508, uc_509, uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, 
      uc_517, uc_518, uc_519, uc_520, uc_521, \P[5] [15], \P[5] [14], \P[5] [13], 
      \P[5] [12], \P[5] [11], \P[5] [10], \P[5] [9], \P[5] [8], \P[5] [7], 
      \P[5] [6], \P[5] [5], \P[5] [4], \P[5] [3], \P[5] [2], \P[5] [1], 
      \P[5] [0], uc_522, uc_523, uc_524, uc_525, uc_526, uc_527, uc_528, uc_529, 
      uc_530, uc_531, uc_532, uc_533, uc_534, uc_535, uc_536, uc_537}), .z({
      uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, uc_546, 
      uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, uc_555, 
      uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, 
      uc_565, uc_566, uc_567, uc_568, \couple[2] [32], \couple[2] [31], 
      \couple[2] [30], \couple[2] [29], \couple[2] [28], \couple[2] [27], 
      \couple[2] [26], \couple[2] [25], \couple[2] [24], \couple[2] [23], 
      \couple[2] [22], \couple[2] [21], \couple[2] [20], \couple[2] [19], 
      \couple[2] [18], \couple[2] [17], \couple[2] [16], uc_569, uc_570, uc_571, 
      uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, uc_580, 
      uc_581, uc_582, uc_583, uc_584}), .C());
   WTM8__1_1898 M6 (.A({a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8]}), 
      .B({b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16]}), .Result(
      \P[6] ));
   WTM8__1_2152 M7 (.A({a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8]}), 
      .B({b[31], b[30], b[29], b[28], b[27], b[26], b[25], b[24]}), .Result(
      \P[7] ));
   adder64__1_3371 A3 (.x({uc_585, uc_586, uc_587, uc_588, uc_589, uc_590, 
      uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, 
      uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, uc_607, uc_608, 
      \P[6] [15], \P[6] [14], \P[6] [13], \P[6] [12], \P[6] [11], \P[6] [10], 
      \P[6] [9], \P[6] [8], uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, 
      uc_615, uc_616, uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, uc_623, 
      uc_624, uc_625, uc_626, uc_627, uc_628, uc_629, uc_630, uc_631, uc_632, 
      uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639, uc_640}), .y({
      uc_641, uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, 
      uc_650, uc_651, uc_652, uc_653, uc_654, uc_655, uc_656, \P[7] [15], 
      \P[7] [14], \P[7] [13], \P[7] [12], \P[7] [11], \P[7] [10], \P[7] [9], 
      \P[7] [8], \P[7] [7], \P[7] [6], \P[7] [5], \P[7] [4], \P[7] [3], 
      \P[7] [2], \P[7] [1], \P[7] [0], uc_657, uc_658, uc_659, uc_660, uc_661, 
      uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, uc_668, uc_669, uc_670, 
      uc_671, uc_672, uc_673, uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, 
      uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, uc_686, uc_687, uc_688}), 
      .z({uc_689, uc_690, uc_691, uc_692, uc_693, uc_694, uc_695, uc_696, uc_697, 
      uc_698, uc_699, uc_700, uc_701, uc_702, uc_703, \couple[3] [48], 
      \couple[3] [47], \couple[3] [46], \couple[3] [45], \couple[3] [44], 
      \couple[3] [43], \couple[3] [42], \couple[3] [41], \couple[3] [40], 
      \couple[3] [39], \couple[3] [38], \couple[3] [37], \couple[3] [36], 
      \couple[3] [35], \couple[3] [34], \couple[3] [33], \couple[3] [32], uc_704, 
      uc_705, uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, uc_712, uc_713, 
      uc_714, uc_715, uc_716, uc_717, uc_718, uc_719, uc_720, uc_721, uc_722, 
      uc_723, uc_724, uc_725, uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, 
      uc_732, uc_733, uc_734, uc_735}), .C());
   adder64__1_3564 A9 (.x({uc_736, uc_737, uc_738, uc_739, uc_740, uc_741, 
      uc_742, uc_743, uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, 
      uc_751, uc_752, uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, 
      uc_760, uc_761, uc_762, uc_763, uc_764, uc_765, uc_766, \couple[2] [32], 
      \couple[2] [31], \couple[2] [30], \couple[2] [29], \couple[2] [28], 
      \couple[2] [27], \couple[2] [26], \couple[2] [25], \couple[2] [24], uc_767, 
      uc_768, uc_769, uc_770, uc_771, uc_772, uc_773, uc_774, uc_775, uc_776, 
      uc_777, uc_778, uc_779, uc_780, uc_781, uc_782, uc_783, uc_784, uc_785, 
      uc_786, uc_787, uc_788, uc_789, uc_790}), .y({uc_791, uc_792, uc_793, 
      uc_794, uc_795, uc_796, uc_797, uc_798, uc_799, uc_800, uc_801, uc_802, 
      uc_803, uc_804, uc_805, \couple[3] [48], \couple[3] [47], \couple[3] [46], 
      \couple[3] [45], \couple[3] [44], \couple[3] [43], \couple[3] [42], 
      \couple[3] [41], \couple[3] [40], \couple[3] [39], \couple[3] [38], 
      \couple[3] [37], \couple[3] [36], \couple[3] [35], \couple[3] [34], 
      \couple[3] [33], \couple[3] [32], \P[6] [7], \P[6] [6], \P[6] [5], 
      \P[6] [4], \P[6] [3], \P[6] [2], \P[6] [1], \P[6] [0], uc_806, uc_807, 
      uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, 
      uc_817, uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, 
      uc_826, uc_827, uc_828, uc_829}), .z({uc_830, uc_831, uc_832, uc_833, 
      uc_834, uc_835, uc_836, uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, 
      uc_843, \Quadruple[1] [49], \Quadruple[1] [48], \Quadruple[1] [47], 
      \Quadruple[1] [46], \Quadruple[1] [45], \Quadruple[1] [44], 
      \Quadruple[1] [43], \Quadruple[1] [42], \Quadruple[1] [41], 
      \Quadruple[1] [40], \Quadruple[1] [39], \Quadruple[1] [38], 
      \Quadruple[1] [37], \Quadruple[1] [36], \Quadruple[1] [35], 
      \Quadruple[1] [34], \Quadruple[1] [33], \Quadruple[1] [32], 
      \Quadruple[1] [31], \Quadruple[1] [30], \Quadruple[1] [29], 
      \Quadruple[1] [28], \Quadruple[1] [27], \Quadruple[1] [26], 
      \Quadruple[1] [25], \Quadruple[1] [24], uc_844, uc_845, uc_846, uc_847, 
      uc_848, uc_849, uc_850, uc_851, uc_852, uc_853, uc_854, uc_855, uc_856, 
      uc_857, uc_858, uc_859, uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, 
      uc_866, uc_867}), .C());
   adder64__1_3757 A12 (.x({uc_868, uc_869, uc_870, uc_871, uc_872, uc_873, 
      uc_874, uc_875, uc_876, uc_877, uc_878, uc_879, uc_880, uc_881, uc_882, 
      uc_883, uc_884, uc_885, uc_886, uc_887, uc_888, uc_889, \Quadruple[0] [41], 
      \Quadruple[0] [40], \Quadruple[0] [39], \Quadruple[0] [38], 
      \Quadruple[0] [37], \Quadruple[0] [36], \Quadruple[0] [35], 
      \Quadruple[0] [34], \Quadruple[0] [33], \Quadruple[0] [32], 
      \Quadruple[0] [31], \Quadruple[0] [30], \Quadruple[0] [29], 
      \Quadruple[0] [28], \Quadruple[0] [27], \Quadruple[0] [26], 
      \Quadruple[0] [25], \Quadruple[0] [24], \Quadruple[0] [23], 
      \Quadruple[0] [22], \Quadruple[0] [21], \Quadruple[0] [20], 
      \Quadruple[0] [19], \Quadruple[0] [18], \Quadruple[0] [17], 
      \Quadruple[0] [16], \couple[0] [15], \couple[0] [14], \couple[0] [13], 
      \couple[0] [12], \couple[0] [11], \couple[0] [10], \couple[0] [9], 
      \couple[0] [8], uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, uc_896, 
      uc_897}), .y({uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, 
      uc_905, uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, \Quadruple[1] [49], 
      \Quadruple[1] [48], \Quadruple[1] [47], \Quadruple[1] [46], 
      \Quadruple[1] [45], \Quadruple[1] [44], \Quadruple[1] [43], 
      \Quadruple[1] [42], \Quadruple[1] [41], \Quadruple[1] [40], 
      \Quadruple[1] [39], \Quadruple[1] [38], \Quadruple[1] [37], 
      \Quadruple[1] [36], \Quadruple[1] [35], \Quadruple[1] [34], 
      \Quadruple[1] [33], \Quadruple[1] [32], \Quadruple[1] [31], 
      \Quadruple[1] [30], \Quadruple[1] [29], \Quadruple[1] [28], 
      \Quadruple[1] [27], \Quadruple[1] [26], \Quadruple[1] [25], 
      \Quadruple[1] [24], \couple[2] [23], \couple[2] [22], \couple[2] [21], 
      \couple[2] [20], \couple[2] [19], \couple[2] [18], \couple[2] [17], 
      \couple[2] [16], \P[4] [7], \P[4] [6], \P[4] [5], \P[4] [4], \P[4] [3], 
      \P[4] [2], \P[4] [1], \P[4] [0], uc_912, uc_913, uc_914, uc_915, uc_916, 
      uc_917, uc_918, uc_919}), .z({uc_920, uc_921, uc_922, uc_923, uc_924, 
      uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, 
      \Eight[0] [50], \Eight[0] [49], \Eight[0] [48], \Eight[0] [47], 
      \Eight[0] [46], \Eight[0] [45], \Eight[0] [44], \Eight[0] [43], 
      \Eight[0] [42], \Eight[0] [41], \Eight[0] [40], \Eight[0] [39], 
      \Eight[0] [38], \Eight[0] [37], \Eight[0] [36], \Eight[0] [35], 
      \Eight[0] [34], \Eight[0] [33], \Eight[0] [32], \Eight[0] [31], 
      \Eight[0] [30], \Eight[0] [29], \Eight[0] [28], \Eight[0] [27], 
      \Eight[0] [26], \Eight[0] [25], \Eight[0] [24], \Eight[0] [23], 
      \Eight[0] [22], \Eight[0] [21], \Eight[0] [20], \Eight[0] [19], 
      \Eight[0] [18], \Eight[0] [17], \Eight[0] [16], \Eight[0] [15], 
      \Eight[0] [14], \Eight[0] [13], \Eight[0] [12], \Eight[0] [11], 
      \Eight[0] [10], \Eight[0] [9], \Eight[0] [8], uc_933, uc_934, uc_935, 
      uc_936, uc_937, uc_938, uc_939, uc_940}), .C());
   datapath__0_81 i_0_1 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_941}), .B(B));
   datapath__0_79 i_0_3 (.p_0({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
      n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, 
      n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, 
      n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, uc_942}), .A(A));
   WTM8__1_2406 M10 (.A({a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16]}), 
      .B({b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16]}), .Result(
      \P[10] ));
   datapath i_0_6 (.p_0({n_0_62, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, 
      n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
      n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, uc_943}), .out({out[63], out[62], 
      out[61], out[60], out[59], out[58], out[57], out[56], out[55], out[54], 
      out[53], out[52], out[51], out[50], out[49], out[48], out[47], out[46], 
      out[45], out[44], out[43], out[42], out[41], out[40], out[39], out[38], 
      out[37], out[36], out[35], out[34], out[33], out[32], out[31], out[30], 
      out[29], out[28], out[27], out[26], out[25], out[24], out[23], out[22], 
      out[21], out[20], out[19], out[18], out[17], out[16], \Eight[0] [15], 
      \Eight[0] [14], \Eight[0] [13], \Eight[0] [12], \Eight[0] [11], 
      \Eight[0] [10], \Eight[0] [9], \Eight[0] [8], \P[0] [7], \P[0] [6], 
      \P[0] [5], \P[0] [4], \P[0] [3], \P[0] [2], \P[0] [1], Result[0]}));
   adder64__0_154 A14 (.x({uc_944, uc_945, uc_946, uc_947, uc_948, uc_949, 
      uc_950, uc_951, uc_952, uc_953, uc_954, uc_955, uc_956, \Eight[0] [50], 
      \Eight[0] [49], \Eight[0] [48], \Eight[0] [47], \Eight[0] [46], 
      \Eight[0] [45], \Eight[0] [44], \Eight[0] [43], \Eight[0] [42], 
      \Eight[0] [41], \Eight[0] [40], \Eight[0] [39], \Eight[0] [38], 
      \Eight[0] [37], \Eight[0] [36], \Eight[0] [35], \Eight[0] [34], 
      \Eight[0] [33], \Eight[0] [32], \Eight[0] [31], \Eight[0] [30], 
      \Eight[0] [29], \Eight[0] [28], \Eight[0] [27], \Eight[0] [26], 
      \Eight[0] [25], \Eight[0] [24], \Eight[0] [23], \Eight[0] [22], 
      \Eight[0] [21], \Eight[0] [20], \Eight[0] [19], \Eight[0] [18], 
      \Eight[0] [17], \Eight[0] [16], uc_957, uc_958, uc_959, uc_960, uc_961, 
      uc_962, uc_963, uc_964, uc_965, uc_966, uc_967, uc_968, uc_969, uc_970, 
      uc_971, uc_972}), .y({\Eight[1] [63], \Eight[1] [62], \Eight[1] [61], 
      \Eight[1] [60], \Eight[1] [59], \Eight[1] [58], \Eight[1] [57], 
      \Eight[1] [56], \Eight[1] [55], \Eight[1] [54], \Eight[1] [53], 
      \Eight[1] [52], \Eight[1] [51], \Eight[1] [50], \Eight[1] [49], 
      \Eight[1] [48], \Eight[1] [47], \Eight[1] [46], \Eight[1] [45], 
      \Eight[1] [44], \Eight[1] [43], \Eight[1] [42], \Eight[1] [41], 
      \Eight[1] [40], \Eight[1] [39], \Eight[1] [38], \Eight[1] [37], 
      \Eight[1] [36], \Eight[1] [35], \Eight[1] [34], \Eight[1] [33], 
      \Eight[1] [32], \Eight[1] [31], \Eight[1] [30], \Eight[1] [29], 
      \Eight[1] [28], \Eight[1] [27], \Eight[1] [26], \Eight[1] [25], 
      \Eight[1] [24], \Eight[1] [23], \Eight[1] [22], \Eight[1] [21], 
      \Eight[1] [20], \Eight[1] [19], \Eight[1] [18], \Eight[1] [17], 
      \Eight[1] [16], uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, 
      uc_980, uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, uc_987, uc_988}), 
      .z({out[63], out[62], out[61], out[60], out[59], out[58], out[57], out[56], 
      out[55], out[54], out[53], out[52], out[51], out[50], out[49], out[48], 
      out[47], out[46], out[45], out[44], out[43], out[42], out[41], out[40], 
      out[39], out[38], out[37], out[36], out[35], out[34], out[33], out[32], 
      out[31], out[30], out[29], out[28], out[27], out[26], out[25], out[24], 
      out[23], out[22], out[21], out[20], out[19], out[18], out[17], out[16], 
      uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, uc_997, 
      uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004}), .C());
   WTM8__0_153 M14 (.A({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24]}), 
      .B({b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16]}), .Result(
      \P[14] ));
   MUX2_X1 i_0_0_0 (.A(B[1]), .B(n_0_0), .S(B[31]), .Z(b[1]));
   MUX2_X1 i_0_0_1 (.A(B[2]), .B(n_0_1), .S(B[31]), .Z(b[2]));
   MUX2_X1 i_0_0_2 (.A(B[3]), .B(n_0_2), .S(B[31]), .Z(b[3]));
   MUX2_X1 i_0_0_3 (.A(B[4]), .B(n_0_3), .S(B[31]), .Z(b[4]));
   MUX2_X1 i_0_0_4 (.A(B[5]), .B(n_0_4), .S(B[31]), .Z(b[5]));
   MUX2_X1 i_0_0_5 (.A(B[6]), .B(n_0_5), .S(B[31]), .Z(b[6]));
   MUX2_X1 i_0_0_6 (.A(B[7]), .B(n_0_6), .S(B[31]), .Z(b[7]));
   MUX2_X1 i_0_0_7 (.A(B[8]), .B(n_0_7), .S(B[31]), .Z(b[8]));
   MUX2_X1 i_0_0_8 (.A(B[9]), .B(n_0_8), .S(B[31]), .Z(b[9]));
   MUX2_X1 i_0_0_9 (.A(B[10]), .B(n_0_9), .S(B[31]), .Z(b[10]));
   MUX2_X1 i_0_0_10 (.A(B[11]), .B(n_0_10), .S(B[31]), .Z(b[11]));
   MUX2_X1 i_0_0_11 (.A(B[12]), .B(n_0_11), .S(B[31]), .Z(b[12]));
   MUX2_X1 i_0_0_12 (.A(B[13]), .B(n_0_12), .S(B[31]), .Z(b[13]));
   MUX2_X1 i_0_0_13 (.A(B[14]), .B(n_0_13), .S(B[31]), .Z(b[14]));
   MUX2_X1 i_0_0_14 (.A(B[15]), .B(n_0_14), .S(B[31]), .Z(b[15]));
   MUX2_X1 i_0_0_15 (.A(B[16]), .B(n_0_15), .S(B[31]), .Z(b[16]));
   MUX2_X1 i_0_0_16 (.A(B[17]), .B(n_0_16), .S(B[31]), .Z(b[17]));
   MUX2_X1 i_0_0_17 (.A(B[18]), .B(n_0_17), .S(B[31]), .Z(b[18]));
   MUX2_X1 i_0_0_18 (.A(B[19]), .B(n_0_18), .S(B[31]), .Z(b[19]));
   MUX2_X1 i_0_0_19 (.A(B[20]), .B(n_0_19), .S(B[31]), .Z(b[20]));
   MUX2_X1 i_0_0_20 (.A(B[21]), .B(n_0_20), .S(B[31]), .Z(b[21]));
   MUX2_X1 i_0_0_21 (.A(B[22]), .B(n_0_21), .S(B[31]), .Z(b[22]));
   MUX2_X1 i_0_0_22 (.A(B[23]), .B(n_0_22), .S(B[31]), .Z(b[23]));
   MUX2_X1 i_0_0_23 (.A(B[24]), .B(n_0_23), .S(B[31]), .Z(b[24]));
   MUX2_X1 i_0_0_24 (.A(B[25]), .B(n_0_24), .S(B[31]), .Z(b[25]));
   MUX2_X1 i_0_0_25 (.A(B[26]), .B(n_0_25), .S(B[31]), .Z(b[26]));
   MUX2_X1 i_0_0_26 (.A(B[27]), .B(n_0_26), .S(B[31]), .Z(b[27]));
   MUX2_X1 i_0_0_27 (.A(B[28]), .B(n_0_27), .S(B[31]), .Z(b[28]));
   MUX2_X1 i_0_0_28 (.A(B[29]), .B(n_0_28), .S(B[31]), .Z(b[29]));
   MUX2_X1 i_0_0_29 (.A(B[30]), .B(n_0_29), .S(B[31]), .Z(b[30]));
   AND2_X1 i_0_0_30 (.A1(n_0_30), .A2(B[31]), .ZN(b[31]));
   MUX2_X1 i_0_0_31 (.A(A[1]), .B(n_0_31), .S(A[31]), .Z(a[1]));
   MUX2_X1 i_0_0_32 (.A(A[2]), .B(n_0_32), .S(A[31]), .Z(a[2]));
   MUX2_X1 i_0_0_33 (.A(A[3]), .B(n_0_33), .S(A[31]), .Z(a[3]));
   MUX2_X1 i_0_0_34 (.A(A[4]), .B(n_0_34), .S(A[31]), .Z(a[4]));
   MUX2_X1 i_0_0_35 (.A(A[5]), .B(n_0_35), .S(A[31]), .Z(a[5]));
   MUX2_X1 i_0_0_36 (.A(A[6]), .B(n_0_36), .S(A[31]), .Z(a[6]));
   MUX2_X1 i_0_0_37 (.A(A[7]), .B(n_0_37), .S(A[31]), .Z(a[7]));
   MUX2_X1 i_0_0_38 (.A(A[8]), .B(n_0_38), .S(A[31]), .Z(a[8]));
   MUX2_X1 i_0_0_39 (.A(A[9]), .B(n_0_39), .S(A[31]), .Z(a[9]));
   MUX2_X1 i_0_0_40 (.A(A[10]), .B(n_0_40), .S(A[31]), .Z(a[10]));
   MUX2_X1 i_0_0_41 (.A(A[11]), .B(n_0_41), .S(A[31]), .Z(a[11]));
   MUX2_X1 i_0_0_42 (.A(A[12]), .B(n_0_42), .S(A[31]), .Z(a[12]));
   MUX2_X1 i_0_0_43 (.A(A[13]), .B(n_0_43), .S(A[31]), .Z(a[13]));
   MUX2_X1 i_0_0_44 (.A(A[14]), .B(n_0_44), .S(A[31]), .Z(a[14]));
   MUX2_X1 i_0_0_45 (.A(A[15]), .B(n_0_45), .S(A[31]), .Z(a[15]));
   MUX2_X1 i_0_0_46 (.A(A[16]), .B(n_0_46), .S(A[31]), .Z(a[16]));
   MUX2_X1 i_0_0_47 (.A(A[17]), .B(n_0_47), .S(A[31]), .Z(a[17]));
   MUX2_X1 i_0_0_48 (.A(A[18]), .B(n_0_48), .S(A[31]), .Z(a[18]));
   MUX2_X1 i_0_0_49 (.A(A[19]), .B(n_0_49), .S(A[31]), .Z(a[19]));
   MUX2_X1 i_0_0_50 (.A(A[20]), .B(n_0_50), .S(A[31]), .Z(a[20]));
   MUX2_X1 i_0_0_51 (.A(A[21]), .B(n_0_51), .S(A[31]), .Z(a[21]));
   MUX2_X1 i_0_0_52 (.A(A[22]), .B(n_0_52), .S(A[31]), .Z(a[22]));
   MUX2_X1 i_0_0_53 (.A(A[23]), .B(n_0_53), .S(A[31]), .Z(a[23]));
   MUX2_X1 i_0_0_54 (.A(A[24]), .B(n_0_54), .S(A[31]), .Z(a[24]));
   MUX2_X1 i_0_0_55 (.A(A[25]), .B(n_0_55), .S(A[31]), .Z(a[25]));
   MUX2_X1 i_0_0_56 (.A(A[26]), .B(n_0_56), .S(A[31]), .Z(a[26]));
   MUX2_X1 i_0_0_57 (.A(A[27]), .B(n_0_57), .S(A[31]), .Z(a[27]));
   MUX2_X1 i_0_0_58 (.A(A[28]), .B(n_0_58), .S(A[31]), .Z(a[28]));
   MUX2_X1 i_0_0_59 (.A(A[29]), .B(n_0_59), .S(A[31]), .Z(a[29]));
   MUX2_X1 i_0_0_60 (.A(A[30]), .B(n_0_60), .S(A[31]), .Z(a[30]));
   AND2_X1 i_0_0_61 (.A1(n_0_61), .A2(A[31]), .ZN(a[31]));
   XNOR2_X1 i_0_0_62 (.A(B[31]), .B(A[31]), .ZN(n_0_0_0));
   MUX2_X1 i_0_0_63 (.A(n_0_63), .B(\P[0] [1]), .S(n_0_0_0), .Z(Result[1]));
   MUX2_X1 i_0_0_64 (.A(n_0_64), .B(\P[0] [2]), .S(n_0_0_0), .Z(Result[2]));
   MUX2_X1 i_0_0_65 (.A(n_0_65), .B(\P[0] [3]), .S(n_0_0_0), .Z(Result[3]));
   MUX2_X1 i_0_0_66 (.A(n_0_66), .B(\P[0] [4]), .S(n_0_0_0), .Z(Result[4]));
   MUX2_X1 i_0_0_67 (.A(n_0_67), .B(\P[0] [5]), .S(n_0_0_0), .Z(Result[5]));
   MUX2_X1 i_0_0_68 (.A(n_0_68), .B(\P[0] [6]), .S(n_0_0_0), .Z(Result[6]));
   MUX2_X1 i_0_0_69 (.A(n_0_69), .B(\P[0] [7]), .S(n_0_0_0), .Z(Result[7]));
   MUX2_X1 i_0_0_70 (.A(n_0_70), .B(\Eight[0] [8]), .S(n_0_0_0), .Z(Result[8]));
   MUX2_X1 i_0_0_71 (.A(n_0_71), .B(\Eight[0] [9]), .S(n_0_0_0), .Z(Result[9]));
   MUX2_X1 i_0_0_72 (.A(n_0_72), .B(\Eight[0] [10]), .S(n_0_0_0), .Z(Result[10]));
   MUX2_X1 i_0_0_73 (.A(n_0_73), .B(\Eight[0] [11]), .S(n_0_0_0), .Z(Result[11]));
   MUX2_X1 i_0_0_74 (.A(n_0_74), .B(\Eight[0] [12]), .S(n_0_0_0), .Z(Result[12]));
   MUX2_X1 i_0_0_75 (.A(n_0_75), .B(\Eight[0] [13]), .S(n_0_0_0), .Z(Result[13]));
   MUX2_X1 i_0_0_76 (.A(n_0_76), .B(\Eight[0] [14]), .S(n_0_0_0), .Z(Result[14]));
   MUX2_X1 i_0_0_77 (.A(n_0_77), .B(\Eight[0] [15]), .S(n_0_0_0), .Z(Result[15]));
   MUX2_X1 i_0_0_78 (.A(n_0_78), .B(out[16]), .S(n_0_0_0), .Z(Result[16]));
   MUX2_X1 i_0_0_79 (.A(n_0_79), .B(out[17]), .S(n_0_0_0), .Z(Result[17]));
   MUX2_X1 i_0_0_80 (.A(n_0_80), .B(out[18]), .S(n_0_0_0), .Z(Result[18]));
   MUX2_X1 i_0_0_81 (.A(n_0_81), .B(out[19]), .S(n_0_0_0), .Z(Result[19]));
   MUX2_X1 i_0_0_82 (.A(n_0_82), .B(out[20]), .S(n_0_0_0), .Z(Result[20]));
   MUX2_X1 i_0_0_83 (.A(n_0_83), .B(out[21]), .S(n_0_0_0), .Z(Result[21]));
   MUX2_X1 i_0_0_84 (.A(n_0_84), .B(out[22]), .S(n_0_0_0), .Z(Result[22]));
   MUX2_X1 i_0_0_85 (.A(n_0_85), .B(out[23]), .S(n_0_0_0), .Z(Result[23]));
   MUX2_X1 i_0_0_86 (.A(n_0_86), .B(out[24]), .S(n_0_0_0), .Z(Result[24]));
   MUX2_X1 i_0_0_87 (.A(n_0_87), .B(out[25]), .S(n_0_0_0), .Z(Result[25]));
   MUX2_X1 i_0_0_88 (.A(n_0_88), .B(out[26]), .S(n_0_0_0), .Z(Result[26]));
   MUX2_X1 i_0_0_89 (.A(n_0_89), .B(out[27]), .S(n_0_0_0), .Z(Result[27]));
   MUX2_X1 i_0_0_90 (.A(n_0_90), .B(out[28]), .S(n_0_0_0), .Z(Result[28]));
   MUX2_X1 i_0_0_91 (.A(n_0_91), .B(out[29]), .S(n_0_0_0), .Z(Result[29]));
   MUX2_X1 i_0_0_92 (.A(n_0_92), .B(out[30]), .S(n_0_0_0), .Z(Result[30]));
   MUX2_X1 i_0_0_93 (.A(n_0_93), .B(out[31]), .S(n_0_0_0), .Z(Result[31]));
   MUX2_X1 i_0_0_94 (.A(n_0_94), .B(out[32]), .S(n_0_0_0), .Z(Result[32]));
   MUX2_X1 i_0_0_95 (.A(n_0_95), .B(out[33]), .S(n_0_0_0), .Z(Result[33]));
   MUX2_X1 i_0_0_96 (.A(n_0_96), .B(out[34]), .S(n_0_0_0), .Z(Result[34]));
   MUX2_X1 i_0_0_97 (.A(n_0_97), .B(out[35]), .S(n_0_0_0), .Z(Result[35]));
   MUX2_X1 i_0_0_98 (.A(n_0_98), .B(out[36]), .S(n_0_0_0), .Z(Result[36]));
   MUX2_X1 i_0_0_99 (.A(n_0_99), .B(out[37]), .S(n_0_0_0), .Z(Result[37]));
   MUX2_X1 i_0_0_100 (.A(n_0_100), .B(out[38]), .S(n_0_0_0), .Z(Result[38]));
   MUX2_X1 i_0_0_101 (.A(n_0_101), .B(out[39]), .S(n_0_0_0), .Z(Result[39]));
   MUX2_X1 i_0_0_102 (.A(n_0_102), .B(out[40]), .S(n_0_0_0), .Z(Result[40]));
   MUX2_X1 i_0_0_103 (.A(n_0_103), .B(out[41]), .S(n_0_0_0), .Z(Result[41]));
   MUX2_X1 i_0_0_104 (.A(n_0_104), .B(out[42]), .S(n_0_0_0), .Z(Result[42]));
   MUX2_X1 i_0_0_105 (.A(n_0_105), .B(out[43]), .S(n_0_0_0), .Z(Result[43]));
   MUX2_X1 i_0_0_106 (.A(n_0_106), .B(out[44]), .S(n_0_0_0), .Z(Result[44]));
   MUX2_X1 i_0_0_107 (.A(n_0_107), .B(out[45]), .S(n_0_0_0), .Z(Result[45]));
   MUX2_X1 i_0_0_108 (.A(n_0_108), .B(out[46]), .S(n_0_0_0), .Z(Result[46]));
   MUX2_X1 i_0_0_109 (.A(n_0_109), .B(out[47]), .S(n_0_0_0), .Z(Result[47]));
   MUX2_X1 i_0_0_110 (.A(n_0_110), .B(out[48]), .S(n_0_0_0), .Z(Result[48]));
   MUX2_X1 i_0_0_111 (.A(n_0_111), .B(out[49]), .S(n_0_0_0), .Z(Result[49]));
   MUX2_X1 i_0_0_112 (.A(n_0_112), .B(out[50]), .S(n_0_0_0), .Z(Result[50]));
   MUX2_X1 i_0_0_113 (.A(n_0_113), .B(out[51]), .S(n_0_0_0), .Z(Result[51]));
   MUX2_X1 i_0_0_114 (.A(n_0_114), .B(out[52]), .S(n_0_0_0), .Z(Result[52]));
   MUX2_X1 i_0_0_115 (.A(n_0_115), .B(out[53]), .S(n_0_0_0), .Z(Result[53]));
   MUX2_X1 i_0_0_116 (.A(n_0_116), .B(out[54]), .S(n_0_0_0), .Z(Result[54]));
   MUX2_X1 i_0_0_117 (.A(n_0_117), .B(out[55]), .S(n_0_0_0), .Z(Result[55]));
   MUX2_X1 i_0_0_118 (.A(n_0_118), .B(out[56]), .S(n_0_0_0), .Z(Result[56]));
   MUX2_X1 i_0_0_119 (.A(n_0_119), .B(out[57]), .S(n_0_0_0), .Z(Result[57]));
   MUX2_X1 i_0_0_120 (.A(n_0_120), .B(out[58]), .S(n_0_0_0), .Z(Result[58]));
   MUX2_X1 i_0_0_121 (.A(n_0_121), .B(out[59]), .S(n_0_0_0), .Z(Result[59]));
   MUX2_X1 i_0_0_122 (.A(n_0_122), .B(out[60]), .S(n_0_0_0), .Z(Result[60]));
   MUX2_X1 i_0_0_123 (.A(n_0_123), .B(out[61]), .S(n_0_0_0), .Z(Result[61]));
   MUX2_X1 i_0_0_124 (.A(n_0_124), .B(out[62]), .S(n_0_0_0), .Z(Result[62]));
   MUX2_X1 i_0_0_125 (.A(n_0_62), .B(out[63]), .S(n_0_0_0), .Z(Result[63]));
   adder64__2_2091 A6 (.x({uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, 
      uc_1011, uc_1012, uc_1013, uc_1014, uc_1015, uc_1016, uc_1017, uc_1018, 
      uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, uc_1026, 
      uc_1027, uc_1028, \P[12] [15], \P[12] [14], \P[12] [13], \P[12] [12], 
      \P[12] [11], \P[12] [10], \P[12] [9], \P[12] [8], uc_1029, uc_1030, 
      uc_1031, uc_1032, uc_1033, uc_1034, uc_1035, uc_1036, uc_1037, uc_1038, 
      uc_1039, uc_1040, uc_1041, uc_1042, uc_1043, uc_1044, uc_1045, uc_1046, 
      uc_1047, uc_1048, uc_1049, uc_1050, uc_1051, uc_1052, uc_1053, uc_1054, 
      uc_1055, uc_1056, uc_1057, uc_1058, uc_1059, uc_1060}), .y({uc_1061, 
      uc_1062, uc_1063, uc_1064, uc_1065, uc_1066, uc_1067, uc_1068, uc_1069, 
      uc_1070, uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, uc_1076, \P[13] [15], 
      \P[13] [14], \P[13] [13], \P[13] [12], \P[13] [11], \P[13] [10], 
      \P[13] [9], \P[13] [8], \P[13] [7], \P[13] [6], \P[13] [5], \P[13] [4], 
      \P[13] [3], \P[13] [2], \P[13] [1], \P[13] [0], uc_1077, uc_1078, uc_1079, 
      uc_1080, uc_1081, uc_1082, uc_1083, uc_1084, uc_1085, uc_1086, uc_1087, 
      uc_1088, uc_1089, uc_1090, uc_1091, uc_1092, uc_1093, uc_1094, uc_1095, 
      uc_1096, uc_1097, uc_1098, uc_1099, uc_1100, uc_1101, uc_1102, uc_1103, 
      uc_1104, uc_1105, uc_1106, uc_1107, uc_1108}), .z({uc_1109, uc_1110, 
      uc_1111, uc_1112, uc_1113, uc_1114, uc_1115, uc_1116, uc_1117, uc_1118, 
      uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, \couple[6] [48], 
      \couple[6] [47], \couple[6] [46], \couple[6] [45], \couple[6] [44], 
      \couple[6] [43], \couple[6] [42], \couple[6] [41], \couple[6] [40], 
      \couple[6] [39], \couple[6] [38], \couple[6] [37], \couple[6] [36], 
      \couple[6] [35], \couple[6] [34], \couple[6] [33], \couple[6] [32], 
      uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, uc_1131, 
      uc_1132, uc_1133, uc_1134, uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, 
      uc_1140, uc_1141, uc_1142, uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, 
      uc_1148, uc_1149, uc_1150, uc_1151, uc_1152, uc_1153, uc_1154, uc_1155}), 
      .C());
   WTM8__2_628 M13 (.A({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24]}), 
      .B({b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8]}), .Result(
      \P[13] ));
   WTM8__2_882 M15 (.A({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24]}), 
      .B({b[31], b[30], b[29], b[28], b[27], b[26], b[25], b[24]}), .Result(
      \P[15] ));
   adder64__2_2284 A7 (.x({uc_1156, uc_1157, uc_1158, uc_1159, uc_1160, uc_1161, 
      uc_1162, uc_1163, \P[14] [15], \P[14] [14], \P[14] [13], \P[14] [12], 
      \P[14] [11], \P[14] [10], \P[14] [9], \P[14] [8], uc_1164, uc_1165, 
      uc_1166, uc_1167, uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, 
      uc_1174, uc_1175, uc_1176, uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, 
      uc_1182, uc_1183, uc_1184, uc_1185, uc_1186, uc_1187, uc_1188, uc_1189, 
      uc_1190, uc_1191, uc_1192, uc_1193, uc_1194, uc_1195, uc_1196, uc_1197, 
      uc_1198, uc_1199, uc_1200, uc_1201, uc_1202, uc_1203, uc_1204, uc_1205, 
      uc_1206, uc_1207, uc_1208, uc_1209, uc_1210, uc_1211}), .y({\P[15] [15], 
      \P[15] [14], \P[15] [13], \P[15] [12], \P[15] [11], \P[15] [10], 
      \P[15] [9], \P[15] [8], \P[15] [7], \P[15] [6], \P[15] [5], \P[15] [4], 
      \P[15] [3], \P[15] [2], \P[15] [1], \P[15] [0], uc_1212, uc_1213, uc_1214, 
      uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, 
      uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, uc_1230, 
      uc_1231, uc_1232, uc_1233, uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, 
      uc_1239, uc_1240, uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, 
      uc_1247, uc_1248, uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, uc_1254, 
      uc_1255, uc_1256, uc_1257, uc_1258, uc_1259}), .z({\couple[7] [63], 
      \couple[7] [62], \couple[7] [61], \couple[7] [60], \couple[7] [59], 
      \couple[7] [58], \couple[7] [57], \couple[7] [56], \couple[7] [55], 
      \couple[7] [54], \couple[7] [53], \couple[7] [52], \couple[7] [51], 
      \couple[7] [50], \couple[7] [49], \couple[7] [48], uc_1260, uc_1261, 
      uc_1262, uc_1263, uc_1264, uc_1265, uc_1266, uc_1267, uc_1268, uc_1269, 
      uc_1270, uc_1271, uc_1272, uc_1273, uc_1274, uc_1275, uc_1276, uc_1277, 
      uc_1278, uc_1279, uc_1280, uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, 
      uc_1286, uc_1287, uc_1288, uc_1289, uc_1290, uc_1291, uc_1292, uc_1293, 
      uc_1294, uc_1295, uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, uc_1301, 
      uc_1302, uc_1303, uc_1304, uc_1305, uc_1306, uc_1307}), .C());
   adder64__2_2477 A11 (.x({uc_1308, uc_1309, uc_1310, uc_1311, uc_1312, uc_1313, 
      uc_1314, uc_1315, uc_1316, uc_1317, uc_1318, uc_1319, uc_1320, uc_1321, 
      uc_1322, \couple[6] [48], \couple[6] [47], \couple[6] [46], 
      \couple[6] [45], \couple[6] [44], \couple[6] [43], \couple[6] [42], 
      \couple[6] [41], \couple[6] [40], uc_1323, uc_1324, uc_1325, uc_1326, 
      uc_1327, uc_1328, uc_1329, uc_1330, uc_1331, uc_1332, uc_1333, uc_1334, 
      uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, 
      uc_1343, uc_1344, uc_1345, uc_1346, uc_1347, uc_1348, uc_1349, uc_1350, 
      uc_1351, uc_1352, uc_1353, uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, 
      uc_1359, uc_1360, uc_1361, uc_1362}), .y({\couple[7] [63], \couple[7] [62], 
      \couple[7] [61], \couple[7] [60], \couple[7] [59], \couple[7] [58], 
      \couple[7] [57], \couple[7] [56], \couple[7] [55], \couple[7] [54], 
      \couple[7] [53], \couple[7] [52], \couple[7] [51], \couple[7] [50], 
      \couple[7] [49], \couple[7] [48], \P[14] [7], \P[14] [6], \P[14] [5], 
      \P[14] [4], \P[14] [3], \P[14] [2], \P[14] [1], \P[14] [0], uc_1363, 
      uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, uc_1371, 
      uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, uc_1378, uc_1379, 
      uc_1380, uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, 
      uc_1388, uc_1389, uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, 
      uc_1396, uc_1397, uc_1398, uc_1399, uc_1400, uc_1401, uc_1402}), .z({
      \Quadruple[3] [63], \Quadruple[3] [62], \Quadruple[3] [61], 
      \Quadruple[3] [60], \Quadruple[3] [59], \Quadruple[3] [58], 
      \Quadruple[3] [57], \Quadruple[3] [56], \Quadruple[3] [55], 
      \Quadruple[3] [54], \Quadruple[3] [53], \Quadruple[3] [52], 
      \Quadruple[3] [51], \Quadruple[3] [50], \Quadruple[3] [49], 
      \Quadruple[3] [48], \Quadruple[3] [47], \Quadruple[3] [46], 
      \Quadruple[3] [45], \Quadruple[3] [44], \Quadruple[3] [43], 
      \Quadruple[3] [42], \Quadruple[3] [41], \Quadruple[3] [40], uc_1403, 
      uc_1404, uc_1405, uc_1406, uc_1407, uc_1408, uc_1409, uc_1410, uc_1411, 
      uc_1412, uc_1413, uc_1414, uc_1415, uc_1416, uc_1417, uc_1418, uc_1419, 
      uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, uc_1427, 
      uc_1428, uc_1429, uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, uc_1435, 
      uc_1436, uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442}), .C());
   adder64__2_2670 A13 (.x({uc_1443, uc_1444, uc_1445, uc_1446, uc_1447, uc_1448, 
      \Quadruple[2] [57], \Quadruple[2] [56], \Quadruple[2] [55], 
      \Quadruple[2] [54], \Quadruple[2] [53], \Quadruple[2] [52], 
      \Quadruple[2] [51], \Quadruple[2] [50], \Quadruple[2] [49], 
      \Quadruple[2] [48], \Quadruple[2] [47], \Quadruple[2] [46], 
      \Quadruple[2] [45], \Quadruple[2] [44], \Quadruple[2] [43], 
      \Quadruple[2] [42], \Quadruple[2] [41], \Quadruple[2] [40], 
      \Quadruple[2] [39], \Quadruple[2] [38], \Quadruple[2] [37], 
      \Quadruple[2] [36], \Quadruple[2] [35], \Quadruple[2] [34], 
      \Quadruple[2] [33], \Quadruple[2] [32], \couple[4] [31], \couple[4] [30], 
      \couple[4] [29], \couple[4] [28], \couple[4] [27], \couple[4] [26], 
      \couple[4] [25], \couple[4] [24], uc_1449, uc_1450, uc_1451, uc_1452, 
      uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, uc_1458, uc_1459, uc_1460, 
      uc_1461, uc_1462, uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, 
      uc_1469, uc_1470, uc_1471, uc_1472}), .y({\Quadruple[3] [63], 
      \Quadruple[3] [62], \Quadruple[3] [61], \Quadruple[3] [60], 
      \Quadruple[3] [59], \Quadruple[3] [58], \Quadruple[3] [57], 
      \Quadruple[3] [56], \Quadruple[3] [55], \Quadruple[3] [54], 
      \Quadruple[3] [53], \Quadruple[3] [52], \Quadruple[3] [51], 
      \Quadruple[3] [50], \Quadruple[3] [49], \Quadruple[3] [48], 
      \Quadruple[3] [47], \Quadruple[3] [46], \Quadruple[3] [45], 
      \Quadruple[3] [44], \Quadruple[3] [43], \Quadruple[3] [42], 
      \Quadruple[3] [41], \Quadruple[3] [40], \couple[6] [39], \couple[6] [38], 
      \couple[6] [37], \couple[6] [36], \couple[6] [35], \couple[6] [34], 
      \couple[6] [33], \couple[6] [32], \P[12] [7], \P[12] [6], \P[12] [5], 
      \P[12] [4], \P[12] [3], \P[12] [2], \P[12] [1], \P[12] [0], uc_1473, 
      uc_1474, uc_1475, uc_1476, uc_1477, uc_1478, uc_1479, uc_1480, uc_1481, 
      uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, uc_1488, uc_1489, 
      uc_1490, uc_1491, uc_1492, uc_1493, uc_1494, uc_1495, uc_1496}), .z({
      \Eight[1] [63], \Eight[1] [62], \Eight[1] [61], \Eight[1] [60], 
      \Eight[1] [59], \Eight[1] [58], \Eight[1] [57], \Eight[1] [56], 
      \Eight[1] [55], \Eight[1] [54], \Eight[1] [53], \Eight[1] [52], 
      \Eight[1] [51], \Eight[1] [50], \Eight[1] [49], \Eight[1] [48], 
      \Eight[1] [47], \Eight[1] [46], \Eight[1] [45], \Eight[1] [44], 
      \Eight[1] [43], \Eight[1] [42], \Eight[1] [41], \Eight[1] [40], 
      \Eight[1] [39], \Eight[1] [38], \Eight[1] [37], \Eight[1] [36], 
      \Eight[1] [35], \Eight[1] [34], \Eight[1] [33], \Eight[1] [32], 
      \Eight[1] [31], \Eight[1] [30], \Eight[1] [29], \Eight[1] [28], 
      \Eight[1] [27], \Eight[1] [26], \Eight[1] [25], \Eight[1] [24], uc_1497, 
      uc_1498, uc_1499, uc_1500, uc_1501, uc_1502, uc_1503, uc_1504, uc_1505, 
      uc_1506, uc_1507, uc_1508, uc_1509, uc_1510, uc_1511, uc_1512, uc_1513, 
      uc_1514, uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, uc_1520}), .C());
   WTM8__2_1136 M12 (.A({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24]}), 
      .B({b[7], b[6], b[5], b[4], b[3], b[2], b[1], B[0]}), .Result(\P[12] ));
   adder64__2_2863 A10 (.x({uc_1521, uc_1522, uc_1523, uc_1524, uc_1525, uc_1526, 
      uc_1527, uc_1528, uc_1529, uc_1530, uc_1531, uc_1532, uc_1533, uc_1534, 
      uc_1535, uc_1536, uc_1537, uc_1538, uc_1539, uc_1540, uc_1541, uc_1542, 
      uc_1543, \couple[4] [40], \couple[4] [39], \couple[4] [38], 
      \couple[4] [37], \couple[4] [36], \couple[4] [35], \couple[4] [34], 
      \couple[4] [33], \couple[4] [32], uc_1544, uc_1545, uc_1546, uc_1547, 
      uc_1548, uc_1549, uc_1550, uc_1551, uc_1552, uc_1553, uc_1554, uc_1555, 
      uc_1556, uc_1557, uc_1558, uc_1559, uc_1560, uc_1561, uc_1562, uc_1563, 
      uc_1564, uc_1565, uc_1566, uc_1567, uc_1568, uc_1569, uc_1570, uc_1571, 
      uc_1572, uc_1573, uc_1574, uc_1575}), .y({uc_1576, uc_1577, uc_1578, 
      uc_1579, uc_1580, uc_1581, uc_1582, \couple[5] [56], \couple[5] [55], 
      \couple[5] [54], \couple[5] [53], \couple[5] [52], \couple[5] [51], 
      \couple[5] [50], \couple[5] [49], \couple[5] [48], \couple[5] [47], 
      \couple[5] [46], \couple[5] [45], \couple[5] [44], \couple[5] [43], 
      \couple[5] [42], \couple[5] [41], \couple[5] [40], \P[10] [7], \P[10] [6], 
      \P[10] [5], \P[10] [4], \P[10] [3], \P[10] [2], \P[10] [1], \P[10] [0], 
      uc_1583, uc_1584, uc_1585, uc_1586, uc_1587, uc_1588, uc_1589, uc_1590, 
      uc_1591, uc_1592, uc_1593, uc_1594, uc_1595, uc_1596, uc_1597, uc_1598, 
      uc_1599, uc_1600, uc_1601, uc_1602, uc_1603, uc_1604, uc_1605, uc_1606, 
      uc_1607, uc_1608, uc_1609, uc_1610, uc_1611, uc_1612, uc_1613, uc_1614}), 
      .z({uc_1615, uc_1616, uc_1617, uc_1618, uc_1619, uc_1620, 
      \Quadruple[2] [57], \Quadruple[2] [56], \Quadruple[2] [55], 
      \Quadruple[2] [54], \Quadruple[2] [53], \Quadruple[2] [52], 
      \Quadruple[2] [51], \Quadruple[2] [50], \Quadruple[2] [49], 
      \Quadruple[2] [48], \Quadruple[2] [47], \Quadruple[2] [46], 
      \Quadruple[2] [45], \Quadruple[2] [44], \Quadruple[2] [43], 
      \Quadruple[2] [42], \Quadruple[2] [41], \Quadruple[2] [40], 
      \Quadruple[2] [39], \Quadruple[2] [38], \Quadruple[2] [37], 
      \Quadruple[2] [36], \Quadruple[2] [35], \Quadruple[2] [34], 
      \Quadruple[2] [33], \Quadruple[2] [32], uc_1621, uc_1622, uc_1623, uc_1624, 
      uc_1625, uc_1626, uc_1627, uc_1628, uc_1629, uc_1630, uc_1631, uc_1632, 
      uc_1633, uc_1634, uc_1635, uc_1636, uc_1637, uc_1638, uc_1639, uc_1640, 
      uc_1641, uc_1642, uc_1643, uc_1644, uc_1645, uc_1646, uc_1647, uc_1648, 
      uc_1649, uc_1650, uc_1651, uc_1652}), .C());
   adder64__2_3056 A5 (.x({uc_1653, uc_1654, uc_1655, uc_1656, uc_1657, uc_1658, 
      uc_1659, uc_1660, uc_1661, uc_1662, uc_1663, uc_1664, uc_1665, uc_1666, 
      uc_1667, uc_1668, \P[10] [15], \P[10] [14], \P[10] [13], \P[10] [12], 
      \P[10] [11], \P[10] [10], \P[10] [9], \P[10] [8], uc_1669, uc_1670, 
      uc_1671, uc_1672, uc_1673, uc_1674, uc_1675, uc_1676, uc_1677, uc_1678, 
      uc_1679, uc_1680, uc_1681, uc_1682, uc_1683, uc_1684, uc_1685, uc_1686, 
      uc_1687, uc_1688, uc_1689, uc_1690, uc_1691, uc_1692, uc_1693, uc_1694, 
      uc_1695, uc_1696, uc_1697, uc_1698, uc_1699, uc_1700, uc_1701, uc_1702, 
      uc_1703, uc_1704, uc_1705, uc_1706, uc_1707, uc_1708}), .y({uc_1709, 
      uc_1710, uc_1711, uc_1712, uc_1713, uc_1714, uc_1715, uc_1716, \P[11] [15], 
      \P[11] [14], \P[11] [13], \P[11] [12], \P[11] [11], \P[11] [10], 
      \P[11] [9], \P[11] [8], \P[11] [7], \P[11] [6], \P[11] [5], \P[11] [4], 
      \P[11] [3], \P[11] [2], \P[11] [1], \P[11] [0], uc_1717, uc_1718, uc_1719, 
      uc_1720, uc_1721, uc_1722, uc_1723, uc_1724, uc_1725, uc_1726, uc_1727, 
      uc_1728, uc_1729, uc_1730, uc_1731, uc_1732, uc_1733, uc_1734, uc_1735, 
      uc_1736, uc_1737, uc_1738, uc_1739, uc_1740, uc_1741, uc_1742, uc_1743, 
      uc_1744, uc_1745, uc_1746, uc_1747, uc_1748, uc_1749, uc_1750, uc_1751, 
      uc_1752, uc_1753, uc_1754, uc_1755, uc_1756}), .z({uc_1757, uc_1758, 
      uc_1759, uc_1760, uc_1761, uc_1762, uc_1763, \couple[5] [56], 
      \couple[5] [55], \couple[5] [54], \couple[5] [53], \couple[5] [52], 
      \couple[5] [51], \couple[5] [50], \couple[5] [49], \couple[5] [48], 
      \couple[5] [47], \couple[5] [46], \couple[5] [45], \couple[5] [44], 
      \couple[5] [43], \couple[5] [42], \couple[5] [41], \couple[5] [40], 
      uc_1764, uc_1765, uc_1766, uc_1767, uc_1768, uc_1769, uc_1770, uc_1771, 
      uc_1772, uc_1773, uc_1774, uc_1775, uc_1776, uc_1777, uc_1778, uc_1779, 
      uc_1780, uc_1781, uc_1782, uc_1783, uc_1784, uc_1785, uc_1786, uc_1787, 
      uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, uc_1793, uc_1794, uc_1795, 
      uc_1796, uc_1797, uc_1798, uc_1799, uc_1800, uc_1801, uc_1802, uc_1803}), 
      .C());
   WTM8__2_1390 M11 (.A({a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16]}), 
      .B({b[31], b[30], b[29], b[28], b[27], b[26], b[25], b[24]}), .Result(
      \P[11] ));
   adder64 A4 (.x({uc_1804, uc_1805, uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, 
      uc_1811, uc_1812, uc_1813, uc_1814, uc_1815, uc_1816, uc_1817, uc_1818, 
      uc_1819, uc_1820, uc_1821, uc_1822, uc_1823, uc_1824, uc_1825, uc_1826, 
      uc_1827, uc_1828, uc_1829, uc_1830, uc_1831, uc_1832, uc_1833, uc_1834, 
      uc_1835, \P[8] [15], \P[8] [14], \P[8] [13], \P[8] [12], \P[8] [11], 
      \P[8] [10], \P[8] [9], \P[8] [8], uc_1836, uc_1837, uc_1838, uc_1839, 
      uc_1840, uc_1841, uc_1842, uc_1843, uc_1844, uc_1845, uc_1846, uc_1847, 
      uc_1848, uc_1849, uc_1850, uc_1851, uc_1852, uc_1853, uc_1854, uc_1855, 
      uc_1856, uc_1857, uc_1858, uc_1859}), .y({uc_1860, uc_1861, uc_1862, 
      uc_1863, uc_1864, uc_1865, uc_1866, uc_1867, uc_1868, uc_1869, uc_1870, 
      uc_1871, uc_1872, uc_1873, uc_1874, uc_1875, uc_1876, uc_1877, uc_1878, 
      uc_1879, uc_1880, uc_1881, uc_1882, uc_1883, \P[9] [15], \P[9] [14], 
      \P[9] [13], \P[9] [12], \P[9] [11], \P[9] [10], \P[9] [9], \P[9] [8], 
      \P[9] [7], \P[9] [6], \P[9] [5], \P[9] [4], \P[9] [3], \P[9] [2], 
      \P[9] [1], \P[9] [0], uc_1884, uc_1885, uc_1886, uc_1887, uc_1888, uc_1889, 
      uc_1890, uc_1891, uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, uc_1897, 
      uc_1898, uc_1899, uc_1900, uc_1901, uc_1902, uc_1903, uc_1904, uc_1905, 
      uc_1906, uc_1907}), .z({uc_1908, uc_1909, uc_1910, uc_1911, uc_1912, 
      uc_1913, uc_1914, uc_1915, uc_1916, uc_1917, uc_1918, uc_1919, uc_1920, 
      uc_1921, uc_1922, uc_1923, uc_1924, uc_1925, uc_1926, uc_1927, uc_1928, 
      uc_1929, uc_1930, \couple[4] [40], \couple[4] [39], \couple[4] [38], 
      \couple[4] [37], \couple[4] [36], \couple[4] [35], \couple[4] [34], 
      \couple[4] [33], \couple[4] [32], \couple[4] [31], \couple[4] [30], 
      \couple[4] [29], \couple[4] [28], \couple[4] [27], \couple[4] [26], 
      \couple[4] [25], \couple[4] [24], uc_1931, uc_1932, uc_1933, uc_1934, 
      uc_1935, uc_1936, uc_1937, uc_1938, uc_1939, uc_1940, uc_1941, uc_1942, 
      uc_1943, uc_1944, uc_1945, uc_1946, uc_1947, uc_1948, uc_1949, uc_1950, 
      uc_1951, uc_1952, uc_1953, uc_1954}), .C());
   WTM8__2_1644 M9 (.A({a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16]}), 
      .B({b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8]}), .Result(\P[9] ));
   WTM8__2_1898 M8 (.A({a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16]}), 
      .B({b[7], b[6], b[5], b[4], b[3], b[2], b[1], B[0]}), .Result({\P[8] [15], 
      \P[8] [14], \P[8] [13], \P[8] [12], \P[8] [11], \P[8] [10], \P[8] [9], 
      \P[8] [8], \Eight[1] [23], \Eight[1] [22], \Eight[1] [21], \Eight[1] [20], 
      \Eight[1] [19], \Eight[1] [18], \Eight[1] [17], \Eight[1] [16]}));
   WTM8 M1 (.A({a[7], a[6], a[5], a[4], a[3], a[2], a[1], A[0]}), .B({b[15], 
      b[14], b[13], b[12], b[11], b[10], b[9], b[8]}), .Result(\P[1] ));
endmodule

module register__3_1(DATA_IN, DATA_OUT, clk, reset);
   input [31:0]DATA_IN;
   output [31:0]DATA_OUT;
   input clk;
   input reset;

   DFF_X1 \DATA_reg[31]  (.D(n_31), .CK(clk), .Q(DATA_OUT[31]), .QN());
   DFF_X1 \DATA_reg[30]  (.D(n_30), .CK(clk), .Q(DATA_OUT[30]), .QN());
   DFF_X1 \DATA_reg[29]  (.D(n_29), .CK(clk), .Q(DATA_OUT[29]), .QN());
   DFF_X1 \DATA_reg[28]  (.D(n_28), .CK(clk), .Q(DATA_OUT[28]), .QN());
   DFF_X1 \DATA_reg[27]  (.D(n_27), .CK(clk), .Q(DATA_OUT[27]), .QN());
   DFF_X1 \DATA_reg[26]  (.D(n_26), .CK(clk), .Q(DATA_OUT[26]), .QN());
   DFF_X1 \DATA_reg[25]  (.D(n_25), .CK(clk), .Q(DATA_OUT[25]), .QN());
   DFF_X1 \DATA_reg[24]  (.D(n_24), .CK(clk), .Q(DATA_OUT[24]), .QN());
   DFF_X1 \DATA_reg[23]  (.D(n_23), .CK(clk), .Q(DATA_OUT[23]), .QN());
   DFF_X1 \DATA_reg[22]  (.D(n_22), .CK(clk), .Q(DATA_OUT[22]), .QN());
   DFF_X1 \DATA_reg[21]  (.D(n_21), .CK(clk), .Q(DATA_OUT[21]), .QN());
   DFF_X1 \DATA_reg[20]  (.D(n_20), .CK(clk), .Q(DATA_OUT[20]), .QN());
   DFF_X1 \DATA_reg[19]  (.D(n_19), .CK(clk), .Q(DATA_OUT[19]), .QN());
   DFF_X1 \DATA_reg[18]  (.D(n_18), .CK(clk), .Q(DATA_OUT[18]), .QN());
   DFF_X1 \DATA_reg[17]  (.D(n_17), .CK(clk), .Q(DATA_OUT[17]), .QN());
   DFF_X1 \DATA_reg[16]  (.D(n_16), .CK(clk), .Q(DATA_OUT[16]), .QN());
   DFF_X1 \DATA_reg[15]  (.D(n_15), .CK(clk), .Q(DATA_OUT[15]), .QN());
   DFF_X1 \DATA_reg[14]  (.D(n_14), .CK(clk), .Q(DATA_OUT[14]), .QN());
   DFF_X1 \DATA_reg[13]  (.D(n_13), .CK(clk), .Q(DATA_OUT[13]), .QN());
   DFF_X1 \DATA_reg[12]  (.D(n_12), .CK(clk), .Q(DATA_OUT[12]), .QN());
   DFF_X1 \DATA_reg[11]  (.D(n_11), .CK(clk), .Q(DATA_OUT[11]), .QN());
   DFF_X1 \DATA_reg[10]  (.D(n_10), .CK(clk), .Q(DATA_OUT[10]), .QN());
   DFF_X1 \DATA_reg[9]  (.D(n_9), .CK(clk), .Q(DATA_OUT[9]), .QN());
   DFF_X1 \DATA_reg[8]  (.D(n_8), .CK(clk), .Q(DATA_OUT[8]), .QN());
   DFF_X1 \DATA_reg[7]  (.D(n_7), .CK(clk), .Q(DATA_OUT[7]), .QN());
   DFF_X1 \DATA_reg[6]  (.D(n_6), .CK(clk), .Q(DATA_OUT[6]), .QN());
   DFF_X1 \DATA_reg[5]  (.D(n_5), .CK(clk), .Q(DATA_OUT[5]), .QN());
   DFF_X1 \DATA_reg[4]  (.D(n_4), .CK(clk), .Q(DATA_OUT[4]), .QN());
   DFF_X1 \DATA_reg[3]  (.D(n_3), .CK(clk), .Q(DATA_OUT[3]), .QN());
   DFF_X1 \DATA_reg[2]  (.D(n_2), .CK(clk), .Q(DATA_OUT[2]), .QN());
   DFF_X1 \DATA_reg[1]  (.D(n_1), .CK(clk), .Q(DATA_OUT[1]), .QN());
   DFF_X1 \DATA_reg[0]  (.D(n_0), .CK(clk), .Q(DATA_OUT[0]), .QN());
   AND2_X1 i_0_0 (.A1(DATA_IN[0]), .A2(reset), .ZN(n_0));
   AND2_X1 i_0_1 (.A1(reset), .A2(DATA_IN[1]), .ZN(n_1));
   AND2_X1 i_0_2 (.A1(reset), .A2(DATA_IN[2]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(reset), .A2(DATA_IN[3]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(reset), .A2(DATA_IN[4]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(reset), .A2(DATA_IN[5]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(reset), .A2(DATA_IN[6]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(reset), .A2(DATA_IN[7]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(reset), .A2(DATA_IN[8]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(reset), .A2(DATA_IN[9]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(reset), .A2(DATA_IN[10]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(reset), .A2(DATA_IN[11]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(reset), .A2(DATA_IN[12]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(reset), .A2(DATA_IN[13]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(reset), .A2(DATA_IN[14]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(reset), .A2(DATA_IN[15]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(reset), .A2(DATA_IN[16]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(reset), .A2(DATA_IN[17]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(reset), .A2(DATA_IN[18]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(reset), .A2(DATA_IN[19]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(reset), .A2(DATA_IN[20]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(reset), .A2(DATA_IN[21]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(reset), .A2(DATA_IN[22]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(reset), .A2(DATA_IN[23]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(reset), .A2(DATA_IN[24]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(reset), .A2(DATA_IN[25]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(reset), .A2(DATA_IN[26]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(reset), .A2(DATA_IN[27]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(reset), .A2(DATA_IN[28]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(reset), .A2(DATA_IN[29]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(reset), .A2(DATA_IN[30]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(reset), .A2(DATA_IN[31]), .ZN(n_31));
endmodule

module register(DATA_IN, DATA_OUT, clk, reset);
   input [31:0]DATA_IN;
   output [31:0]DATA_OUT;
   input clk;
   input reset;

   DFF_X1 \DATA_reg[31]  (.D(n_31), .CK(clk), .Q(DATA_OUT[31]), .QN());
   DFF_X1 \DATA_reg[30]  (.D(n_30), .CK(clk), .Q(DATA_OUT[30]), .QN());
   DFF_X1 \DATA_reg[29]  (.D(n_29), .CK(clk), .Q(DATA_OUT[29]), .QN());
   DFF_X1 \DATA_reg[28]  (.D(n_28), .CK(clk), .Q(DATA_OUT[28]), .QN());
   DFF_X1 \DATA_reg[27]  (.D(n_27), .CK(clk), .Q(DATA_OUT[27]), .QN());
   DFF_X1 \DATA_reg[26]  (.D(n_26), .CK(clk), .Q(DATA_OUT[26]), .QN());
   DFF_X1 \DATA_reg[25]  (.D(n_25), .CK(clk), .Q(DATA_OUT[25]), .QN());
   DFF_X1 \DATA_reg[24]  (.D(n_24), .CK(clk), .Q(DATA_OUT[24]), .QN());
   DFF_X1 \DATA_reg[23]  (.D(n_23), .CK(clk), .Q(DATA_OUT[23]), .QN());
   DFF_X1 \DATA_reg[22]  (.D(n_22), .CK(clk), .Q(DATA_OUT[22]), .QN());
   DFF_X1 \DATA_reg[21]  (.D(n_21), .CK(clk), .Q(DATA_OUT[21]), .QN());
   DFF_X1 \DATA_reg[20]  (.D(n_20), .CK(clk), .Q(DATA_OUT[20]), .QN());
   DFF_X1 \DATA_reg[19]  (.D(n_19), .CK(clk), .Q(DATA_OUT[19]), .QN());
   DFF_X1 \DATA_reg[18]  (.D(n_18), .CK(clk), .Q(DATA_OUT[18]), .QN());
   DFF_X1 \DATA_reg[17]  (.D(n_17), .CK(clk), .Q(DATA_OUT[17]), .QN());
   DFF_X1 \DATA_reg[16]  (.D(n_16), .CK(clk), .Q(DATA_OUT[16]), .QN());
   DFF_X1 \DATA_reg[15]  (.D(n_15), .CK(clk), .Q(DATA_OUT[15]), .QN());
   DFF_X1 \DATA_reg[14]  (.D(n_14), .CK(clk), .Q(DATA_OUT[14]), .QN());
   DFF_X1 \DATA_reg[13]  (.D(n_13), .CK(clk), .Q(DATA_OUT[13]), .QN());
   DFF_X1 \DATA_reg[12]  (.D(n_12), .CK(clk), .Q(DATA_OUT[12]), .QN());
   DFF_X1 \DATA_reg[11]  (.D(n_11), .CK(clk), .Q(DATA_OUT[11]), .QN());
   DFF_X1 \DATA_reg[10]  (.D(n_10), .CK(clk), .Q(DATA_OUT[10]), .QN());
   DFF_X1 \DATA_reg[9]  (.D(n_9), .CK(clk), .Q(DATA_OUT[9]), .QN());
   DFF_X1 \DATA_reg[8]  (.D(n_8), .CK(clk), .Q(DATA_OUT[8]), .QN());
   DFF_X1 \DATA_reg[7]  (.D(n_7), .CK(clk), .Q(DATA_OUT[7]), .QN());
   DFF_X1 \DATA_reg[6]  (.D(n_6), .CK(clk), .Q(DATA_OUT[6]), .QN());
   DFF_X1 \DATA_reg[5]  (.D(n_5), .CK(clk), .Q(DATA_OUT[5]), .QN());
   DFF_X1 \DATA_reg[4]  (.D(n_4), .CK(clk), .Q(DATA_OUT[4]), .QN());
   DFF_X1 \DATA_reg[3]  (.D(n_3), .CK(clk), .Q(DATA_OUT[3]), .QN());
   DFF_X1 \DATA_reg[2]  (.D(n_2), .CK(clk), .Q(DATA_OUT[2]), .QN());
   DFF_X1 \DATA_reg[1]  (.D(n_1), .CK(clk), .Q(DATA_OUT[1]), .QN());
   DFF_X1 \DATA_reg[0]  (.D(n_0), .CK(clk), .Q(DATA_OUT[0]), .QN());
   AND2_X1 i_0_0 (.A1(DATA_IN[0]), .A2(reset), .ZN(n_0));
   AND2_X1 i_0_1 (.A1(reset), .A2(DATA_IN[1]), .ZN(n_1));
   AND2_X1 i_0_2 (.A1(reset), .A2(DATA_IN[2]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(reset), .A2(DATA_IN[3]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(reset), .A2(DATA_IN[4]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(reset), .A2(DATA_IN[5]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(reset), .A2(DATA_IN[6]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(reset), .A2(DATA_IN[7]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(reset), .A2(DATA_IN[8]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(reset), .A2(DATA_IN[9]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(reset), .A2(DATA_IN[10]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(reset), .A2(DATA_IN[11]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(reset), .A2(DATA_IN[12]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(reset), .A2(DATA_IN[13]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(reset), .A2(DATA_IN[14]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(reset), .A2(DATA_IN[15]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(reset), .A2(DATA_IN[16]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(reset), .A2(DATA_IN[17]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(reset), .A2(DATA_IN[18]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(reset), .A2(DATA_IN[19]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(reset), .A2(DATA_IN[20]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(reset), .A2(DATA_IN[21]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(reset), .A2(DATA_IN[22]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(reset), .A2(DATA_IN[23]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(reset), .A2(DATA_IN[24]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(reset), .A2(DATA_IN[25]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(reset), .A2(DATA_IN[26]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(reset), .A2(DATA_IN[27]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(reset), .A2(DATA_IN[28]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(reset), .A2(DATA_IN[29]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(reset), .A2(DATA_IN[30]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(reset), .A2(DATA_IN[31]), .ZN(n_31));
endmodule

module register__parameterized0(DATA_IN, DATA_OUT, clk, reset);
   input [63:0]DATA_IN;
   output [63:0]DATA_OUT;
   input clk;
   input reset;

   DFF_X1 \DATA_reg[63]  (.D(n_63), .CK(clk), .Q(DATA_OUT[63]), .QN());
   DFF_X1 \DATA_reg[62]  (.D(n_62), .CK(clk), .Q(DATA_OUT[62]), .QN());
   DFF_X1 \DATA_reg[61]  (.D(n_61), .CK(clk), .Q(DATA_OUT[61]), .QN());
   DFF_X1 \DATA_reg[60]  (.D(n_60), .CK(clk), .Q(DATA_OUT[60]), .QN());
   DFF_X1 \DATA_reg[59]  (.D(n_59), .CK(clk), .Q(DATA_OUT[59]), .QN());
   DFF_X1 \DATA_reg[58]  (.D(n_58), .CK(clk), .Q(DATA_OUT[58]), .QN());
   DFF_X1 \DATA_reg[57]  (.D(n_57), .CK(clk), .Q(DATA_OUT[57]), .QN());
   DFF_X1 \DATA_reg[56]  (.D(n_56), .CK(clk), .Q(DATA_OUT[56]), .QN());
   DFF_X1 \DATA_reg[55]  (.D(n_55), .CK(clk), .Q(DATA_OUT[55]), .QN());
   DFF_X1 \DATA_reg[54]  (.D(n_54), .CK(clk), .Q(DATA_OUT[54]), .QN());
   DFF_X1 \DATA_reg[53]  (.D(n_53), .CK(clk), .Q(DATA_OUT[53]), .QN());
   DFF_X1 \DATA_reg[52]  (.D(n_52), .CK(clk), .Q(DATA_OUT[52]), .QN());
   DFF_X1 \DATA_reg[51]  (.D(n_51), .CK(clk), .Q(DATA_OUT[51]), .QN());
   DFF_X1 \DATA_reg[50]  (.D(n_50), .CK(clk), .Q(DATA_OUT[50]), .QN());
   DFF_X1 \DATA_reg[49]  (.D(n_49), .CK(clk), .Q(DATA_OUT[49]), .QN());
   DFF_X1 \DATA_reg[48]  (.D(n_48), .CK(clk), .Q(DATA_OUT[48]), .QN());
   DFF_X1 \DATA_reg[47]  (.D(n_47), .CK(clk), .Q(DATA_OUT[47]), .QN());
   DFF_X1 \DATA_reg[46]  (.D(n_46), .CK(clk), .Q(DATA_OUT[46]), .QN());
   DFF_X1 \DATA_reg[45]  (.D(n_45), .CK(clk), .Q(DATA_OUT[45]), .QN());
   DFF_X1 \DATA_reg[44]  (.D(n_44), .CK(clk), .Q(DATA_OUT[44]), .QN());
   DFF_X1 \DATA_reg[43]  (.D(n_43), .CK(clk), .Q(DATA_OUT[43]), .QN());
   DFF_X1 \DATA_reg[42]  (.D(n_42), .CK(clk), .Q(DATA_OUT[42]), .QN());
   DFF_X1 \DATA_reg[41]  (.D(n_41), .CK(clk), .Q(DATA_OUT[41]), .QN());
   DFF_X1 \DATA_reg[40]  (.D(n_40), .CK(clk), .Q(DATA_OUT[40]), .QN());
   DFF_X1 \DATA_reg[39]  (.D(n_39), .CK(clk), .Q(DATA_OUT[39]), .QN());
   DFF_X1 \DATA_reg[38]  (.D(n_38), .CK(clk), .Q(DATA_OUT[38]), .QN());
   DFF_X1 \DATA_reg[37]  (.D(n_37), .CK(clk), .Q(DATA_OUT[37]), .QN());
   DFF_X1 \DATA_reg[36]  (.D(n_36), .CK(clk), .Q(DATA_OUT[36]), .QN());
   DFF_X1 \DATA_reg[35]  (.D(n_35), .CK(clk), .Q(DATA_OUT[35]), .QN());
   DFF_X1 \DATA_reg[34]  (.D(n_34), .CK(clk), .Q(DATA_OUT[34]), .QN());
   DFF_X1 \DATA_reg[33]  (.D(n_33), .CK(clk), .Q(DATA_OUT[33]), .QN());
   DFF_X1 \DATA_reg[32]  (.D(n_32), .CK(clk), .Q(DATA_OUT[32]), .QN());
   DFF_X1 \DATA_reg[31]  (.D(n_31), .CK(clk), .Q(DATA_OUT[31]), .QN());
   DFF_X1 \DATA_reg[30]  (.D(n_30), .CK(clk), .Q(DATA_OUT[30]), .QN());
   DFF_X1 \DATA_reg[29]  (.D(n_29), .CK(clk), .Q(DATA_OUT[29]), .QN());
   DFF_X1 \DATA_reg[28]  (.D(n_28), .CK(clk), .Q(DATA_OUT[28]), .QN());
   DFF_X1 \DATA_reg[27]  (.D(n_27), .CK(clk), .Q(DATA_OUT[27]), .QN());
   DFF_X1 \DATA_reg[26]  (.D(n_26), .CK(clk), .Q(DATA_OUT[26]), .QN());
   DFF_X1 \DATA_reg[25]  (.D(n_25), .CK(clk), .Q(DATA_OUT[25]), .QN());
   DFF_X1 \DATA_reg[24]  (.D(n_24), .CK(clk), .Q(DATA_OUT[24]), .QN());
   DFF_X1 \DATA_reg[23]  (.D(n_23), .CK(clk), .Q(DATA_OUT[23]), .QN());
   DFF_X1 \DATA_reg[22]  (.D(n_22), .CK(clk), .Q(DATA_OUT[22]), .QN());
   DFF_X1 \DATA_reg[21]  (.D(n_21), .CK(clk), .Q(DATA_OUT[21]), .QN());
   DFF_X1 \DATA_reg[20]  (.D(n_20), .CK(clk), .Q(DATA_OUT[20]), .QN());
   DFF_X1 \DATA_reg[19]  (.D(n_19), .CK(clk), .Q(DATA_OUT[19]), .QN());
   DFF_X1 \DATA_reg[18]  (.D(n_18), .CK(clk), .Q(DATA_OUT[18]), .QN());
   DFF_X1 \DATA_reg[17]  (.D(n_17), .CK(clk), .Q(DATA_OUT[17]), .QN());
   DFF_X1 \DATA_reg[16]  (.D(n_16), .CK(clk), .Q(DATA_OUT[16]), .QN());
   DFF_X1 \DATA_reg[15]  (.D(n_15), .CK(clk), .Q(DATA_OUT[15]), .QN());
   DFF_X1 \DATA_reg[14]  (.D(n_14), .CK(clk), .Q(DATA_OUT[14]), .QN());
   DFF_X1 \DATA_reg[13]  (.D(n_13), .CK(clk), .Q(DATA_OUT[13]), .QN());
   DFF_X1 \DATA_reg[12]  (.D(n_12), .CK(clk), .Q(DATA_OUT[12]), .QN());
   DFF_X1 \DATA_reg[11]  (.D(n_11), .CK(clk), .Q(DATA_OUT[11]), .QN());
   DFF_X1 \DATA_reg[10]  (.D(n_10), .CK(clk), .Q(DATA_OUT[10]), .QN());
   DFF_X1 \DATA_reg[9]  (.D(n_9), .CK(clk), .Q(DATA_OUT[9]), .QN());
   DFF_X1 \DATA_reg[8]  (.D(n_8), .CK(clk), .Q(DATA_OUT[8]), .QN());
   DFF_X1 \DATA_reg[7]  (.D(n_7), .CK(clk), .Q(DATA_OUT[7]), .QN());
   DFF_X1 \DATA_reg[6]  (.D(n_6), .CK(clk), .Q(DATA_OUT[6]), .QN());
   DFF_X1 \DATA_reg[5]  (.D(n_5), .CK(clk), .Q(DATA_OUT[5]), .QN());
   DFF_X1 \DATA_reg[4]  (.D(n_4), .CK(clk), .Q(DATA_OUT[4]), .QN());
   DFF_X1 \DATA_reg[3]  (.D(n_3), .CK(clk), .Q(DATA_OUT[3]), .QN());
   DFF_X1 \DATA_reg[2]  (.D(n_2), .CK(clk), .Q(DATA_OUT[2]), .QN());
   DFF_X1 \DATA_reg[1]  (.D(n_1), .CK(clk), .Q(DATA_OUT[1]), .QN());
   DFF_X1 \DATA_reg[0]  (.D(n_0), .CK(clk), .Q(DATA_OUT[0]), .QN());
   AND2_X1 i_0_0 (.A1(DATA_IN[0]), .A2(reset), .ZN(n_0));
   AND2_X1 i_0_1 (.A1(reset), .A2(DATA_IN[1]), .ZN(n_1));
   AND2_X1 i_0_2 (.A1(reset), .A2(DATA_IN[2]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(reset), .A2(DATA_IN[3]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(reset), .A2(DATA_IN[4]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(reset), .A2(DATA_IN[5]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(reset), .A2(DATA_IN[6]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(reset), .A2(DATA_IN[7]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(reset), .A2(DATA_IN[8]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(reset), .A2(DATA_IN[9]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(reset), .A2(DATA_IN[10]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(reset), .A2(DATA_IN[11]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(reset), .A2(DATA_IN[12]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(reset), .A2(DATA_IN[13]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(reset), .A2(DATA_IN[14]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(reset), .A2(DATA_IN[15]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(reset), .A2(DATA_IN[16]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(reset), .A2(DATA_IN[17]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(reset), .A2(DATA_IN[18]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(reset), .A2(DATA_IN[19]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(reset), .A2(DATA_IN[20]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(reset), .A2(DATA_IN[21]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(reset), .A2(DATA_IN[22]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(reset), .A2(DATA_IN[23]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(reset), .A2(DATA_IN[24]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(reset), .A2(DATA_IN[25]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(reset), .A2(DATA_IN[26]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(reset), .A2(DATA_IN[27]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(reset), .A2(DATA_IN[28]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(reset), .A2(DATA_IN[29]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(reset), .A2(DATA_IN[30]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(reset), .A2(DATA_IN[31]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(reset), .A2(DATA_IN[32]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(reset), .A2(DATA_IN[33]), .ZN(n_33));
   AND2_X1 i_0_34 (.A1(reset), .A2(DATA_IN[34]), .ZN(n_34));
   AND2_X1 i_0_35 (.A1(reset), .A2(DATA_IN[35]), .ZN(n_35));
   AND2_X1 i_0_36 (.A1(reset), .A2(DATA_IN[36]), .ZN(n_36));
   AND2_X1 i_0_37 (.A1(reset), .A2(DATA_IN[37]), .ZN(n_37));
   AND2_X1 i_0_38 (.A1(reset), .A2(DATA_IN[38]), .ZN(n_38));
   AND2_X1 i_0_39 (.A1(reset), .A2(DATA_IN[39]), .ZN(n_39));
   AND2_X1 i_0_40 (.A1(reset), .A2(DATA_IN[40]), .ZN(n_40));
   AND2_X1 i_0_41 (.A1(reset), .A2(DATA_IN[41]), .ZN(n_41));
   AND2_X1 i_0_42 (.A1(reset), .A2(DATA_IN[42]), .ZN(n_42));
   AND2_X1 i_0_43 (.A1(reset), .A2(DATA_IN[43]), .ZN(n_43));
   AND2_X1 i_0_44 (.A1(reset), .A2(DATA_IN[44]), .ZN(n_44));
   AND2_X1 i_0_45 (.A1(reset), .A2(DATA_IN[45]), .ZN(n_45));
   AND2_X1 i_0_46 (.A1(reset), .A2(DATA_IN[46]), .ZN(n_46));
   AND2_X1 i_0_47 (.A1(reset), .A2(DATA_IN[47]), .ZN(n_47));
   AND2_X1 i_0_48 (.A1(reset), .A2(DATA_IN[48]), .ZN(n_48));
   AND2_X1 i_0_49 (.A1(reset), .A2(DATA_IN[49]), .ZN(n_49));
   AND2_X1 i_0_50 (.A1(reset), .A2(DATA_IN[50]), .ZN(n_50));
   AND2_X1 i_0_51 (.A1(reset), .A2(DATA_IN[51]), .ZN(n_51));
   AND2_X1 i_0_52 (.A1(reset), .A2(DATA_IN[52]), .ZN(n_52));
   AND2_X1 i_0_53 (.A1(reset), .A2(DATA_IN[53]), .ZN(n_53));
   AND2_X1 i_0_54 (.A1(reset), .A2(DATA_IN[54]), .ZN(n_54));
   AND2_X1 i_0_55 (.A1(reset), .A2(DATA_IN[55]), .ZN(n_55));
   AND2_X1 i_0_56 (.A1(reset), .A2(DATA_IN[56]), .ZN(n_56));
   AND2_X1 i_0_57 (.A1(reset), .A2(DATA_IN[57]), .ZN(n_57));
   AND2_X1 i_0_58 (.A1(reset), .A2(DATA_IN[58]), .ZN(n_58));
   AND2_X1 i_0_59 (.A1(reset), .A2(DATA_IN[59]), .ZN(n_59));
   AND2_X1 i_0_60 (.A1(reset), .A2(DATA_IN[60]), .ZN(n_60));
   AND2_X1 i_0_61 (.A1(reset), .A2(DATA_IN[61]), .ZN(n_61));
   AND2_X1 i_0_62 (.A1(reset), .A2(DATA_IN[62]), .ZN(n_62));
   AND2_X1 i_0_63 (.A1(reset), .A2(DATA_IN[63]), .ZN(n_63));
endmodule

module registered_WTM(A, B, Result, clk, reset);
   input [31:0]A;
   input [31:0]B;
   output [63:0]Result;
   input clk;
   input reset;

   wire [63:0]Result_OUT;
   wire [31:0]A_IN;
   wire [31:0]B_IN;

   WTM32 multiplier (.A(A_IN), .B(B_IN), .Result(Result_OUT));
   register__3_1 inputReg_1 (.DATA_IN(A), .DATA_OUT(A_IN), .clk(clk), .reset(
      reset));
   register inputReg_2 (.DATA_IN(B), .DATA_OUT(B_IN), .clk(clk), .reset(reset));
   register__parameterized0 outputReg (.DATA_IN(Result_OUT), .DATA_OUT(Result), 
      .clk(clk), .reset(reset));
endmodule
