
// 	Wed Jan  4 01:59:07 2023
//	vlsi
//	localhost.localdomain

module datapath__0_15 (p_0, accumulator, p_1);

output [63:0] p_1;
input [63:0] accumulator;
input [63:0] p_0;
wire spw_n22;
wire spw_n8;
wire n_0;
wire n_366;
wire n_1;
wire n_365;
wire n_364;
wire n_2;
wire n_369;
wire n_363;
wire n_3;
wire n_370;
wire n_376;
wire n_372;
wire n_361;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_358;
wire n_349;
wire n_11;
wire n_5;
wire n_359;
wire n_353;
wire n_8;
wire n_356;
wire n_354;
wire n_360;
wire n_351;
wire n_347;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_344;
wire n_335;
wire n_19;
wire n_13;
wire n_345;
wire n_339;
wire n_16;
wire n_342;
wire n_340;
wire n_346;
wire n_337;
wire n_333;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_330;
wire n_321;
wire n_27;
wire n_21;
wire n_331;
wire n_325;
wire n_24;
wire n_328;
wire n_326;
wire n_332;
wire n_323;
wire n_319;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_285;
wire n_275;
wire n_35;
wire n_29;
wire n_284;
wire n_287;
wire n_277;
wire n_32;
wire n_286;
wire n_282;
wire n_279;
wire n_289;
wire n_63;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_313;
wire n_257;
wire n_43;
wire n_37;
wire n_312;
wire n_315;
wire n_259;
wire n_40;
wire n_314;
wire n_318;
wire n_261;
wire n_317;
wire n_61;
wire n_50;
wire n_49;
wire n_46;
wire n_47;
wire n_44;
wire n_296;
wire n_269;
wire n_51;
wire n_45;
wire n_295;
wire n_298;
wire n_271;
wire n_48;
wire n_297;
wire n_293;
wire n_273;
wire n_300;
wire n_59;
wire n_58;
wire n_57;
wire n_54;
wire n_55;
wire n_52;
wire n_305;
wire n_263;
wire n_65;
wire n_53;
wire n_304;
wire n_307;
wire n_266;
wire n_56;
wire n_306;
wire n_302;
wire n_267;
wire n_60;
wire n_268;
wire n_292;
wire n_62;
wire n_256;
wire n_310;
wire n_64;
wire n_274;
wire n_281;
wire n_308;
wire n_377;
wire n_373;
wire n_254;
wire n_72;
wire n_71;
wire n_68;
wire n_69;
wire n_66;
wire n_223;
wire n_213;
wire n_73;
wire n_67;
wire n_222;
wire n_225;
wire n_215;
wire n_70;
wire n_224;
wire n_220;
wire n_217;
wire n_227;
wire n_101;
wire n_80;
wire n_79;
wire n_76;
wire n_77;
wire n_74;
wire n_248;
wire n_206;
wire n_81;
wire n_75;
wire n_247;
wire n_250;
wire n_208;
wire n_78;
wire n_249;
wire n_253;
wire n_210;
wire n_252;
wire n_99;
wire n_88;
wire n_87;
wire n_84;
wire n_85;
wire n_82;
wire n_234;
wire n_192;
wire n_89;
wire n_83;
wire n_233;
wire n_236;
wire n_194;
wire n_86;
wire n_235;
wire n_231;
wire n_196;
wire n_238;
wire n_98;
wire n_97;
wire n_95;
wire n_94;
wire n_91;
wire n_90;
wire n_202;
wire n_242;
wire n_199;
wire n_103;
wire n_92;
wire n_93;
wire n_241;
wire n_200;
wire n_96;
wire n_243;
wire n_203;
wire n_204;
wire n_191;
wire n_230;
wire n_100;
wire n_205;
wire n_245;
wire n_102;
wire n_212;
wire n_219;
wire n_244;
wire n_189;
wire n_110;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_186;
wire n_177;
wire n_111;
wire n_105;
wire n_187;
wire n_181;
wire n_108;
wire n_184;
wire n_182;
wire n_188;
wire n_179;
wire n_175;
wire n_118;
wire n_117;
wire n_114;
wire n_115;
wire n_112;
wire n_164;
wire n_154;
wire n_119;
wire n_113;
wire n_163;
wire n_166;
wire n_156;
wire n_116;
wire n_165;
wire n_161;
wire n_158;
wire n_168;
wire n_128;
wire n_127;
wire n_125;
wire n_124;
wire n_121;
wire n_120;
wire n_149;
wire n_172;
wire n_145;
wire n_129;
wire n_122;
wire n_123;
wire n_171;
wire n_146;
wire n_126;
wire n_173;
wire n_150;
wire n_151;
wire n_153;
wire n_160;
wire n_174;
wire n_143;
wire n_142;
wire n_140;
wire n_136;
wire n_141;
wire n_135;
wire n_131;
wire n_130;
wire n_137;
wire n_139;
wire n_133;
wire n_132;
wire n_134;
wire n_138;
wire n_379;
wire n_375;
wire n_371;
wire n_147;
wire n_144;
wire n_152;
wire n_159;
wire n_378;
wire n_374;
wire n_148;
wire n_170;
wire n_169;
wire n_155;
wire n_167;
wire n_162;
wire n_157;
wire n_176;
wire n_180;
wire n_183;
wire n_178;
wire n_185;
wire n_211;
wire n_190;
wire n_218;
wire n_197;
wire n_239;
wire n_229;
wire n_193;
wire n_237;
wire n_232;
wire n_195;
wire n_198;
wire n_201;
wire n_240;
wire n_207;
wire n_251;
wire n_246;
wire n_209;
wire n_228;
wire n_214;
wire n_226;
wire n_221;
wire n_216;
wire n_262;
wire n_255;
wire n_280;
wire n_290;
wire n_291;
wire n_301;
wire n_258;
wire n_316;
wire n_311;
wire n_260;
wire n_303;
wire n_265;
wire n_309;
wire n_264;
wire n_270;
wire n_299;
wire n_294;
wire n_272;
wire n_276;
wire n_288;
wire n_283;
wire n_278;
wire n_320;
wire n_324;
wire n_327;
wire n_322;
wire n_329;
wire n_334;
wire n_338;
wire n_341;
wire n_336;
wire n_343;
wire n_348;
wire n_352;
wire n_355;
wire n_350;
wire n_357;
wire n_362;
wire n_368;
wire n_367;
wire spw__n10;
wire spw__n11;


INV_X1 i_443 (.ZN (n_379), .A (p_0[61]));
INV_X1 i_442 (.ZN (n_378), .A (p_0[59]));
INV_X1 i_441 (.ZN (n_377), .A (p_0[31]));
INV_X1 i_440 (.ZN (n_376), .A (p_0[3]));
INV_X1 i_439 (.ZN (n_375), .A (accumulator[61]));
INV_X1 i_438 (.ZN (n_374), .A (accumulator[59]));
INV_X1 i_437 (.ZN (n_373), .A (accumulator[31]));
INV_X1 i_436 (.ZN (n_372), .A (accumulator[3]));
NOR2_X1 i_435 (.ZN (n_371), .A1 (p_0[60]), .A2 (accumulator[60]));
NAND2_X1 i_434 (.ZN (n_370), .A1 (n_376), .A2 (n_372));
NAND2_X1 i_433 (.ZN (n_369), .A1 (p_0[2]), .A2 (accumulator[2]));
INV_X1 i_432 (.ZN (n_368), .A (n_369));
NOR2_X1 i_431 (.ZN (n_367), .A1 (p_0[1]), .A2 (spw__n11));
NAND2_X1 i_430 (.ZN (n_366), .A1 (p_0[0]), .A2 (accumulator[0]));
NAND2_X1 i_429 (.ZN (n_365), .A1 (p_0[1]), .A2 (spw__n10));
AOI21_X1 i_428 (.ZN (n_364), .A (n_367), .B1 (n_366), .B2 (n_365));
OAI22_X1 i_427 (.ZN (n_363), .A1 (p_0[2]), .A2 (accumulator[2]), .B1 (n_368), .B2 (n_364));
OAI21_X1 i_426 (.ZN (n_362), .A (n_363), .B1 (n_376), .B2 (n_372));
NAND2_X1 i_425 (.ZN (n_361), .A1 (n_370), .A2 (n_362));
NOR2_X1 i_424 (.ZN (n_360), .A1 (p_0[7]), .A2 (accumulator[7]));
NOR2_X1 i_423 (.ZN (n_359), .A1 (p_0[5]), .A2 (accumulator[5]));
NOR2_X1 i_422 (.ZN (n_358), .A1 (p_0[6]), .A2 (accumulator[6]));
OR3_X1 i_421 (.ZN (n_357), .A1 (n_360), .A2 (n_358), .A3 (n_359));
NOR2_X1 i_420 (.ZN (n_356), .A1 (p_0[4]), .A2 (accumulator[4]));
NOR3_X1 i_419 (.ZN (n_355), .A1 (n_357), .A2 (n_356), .A3 (n_361));
NAND2_X1 i_418 (.ZN (n_354), .A1 (p_0[4]), .A2 (accumulator[4]));
NAND2_X1 i_417 (.ZN (n_353), .A1 (p_0[5]), .A2 (accumulator[5]));
AOI21_X1 i_416 (.ZN (n_352), .A (n_357), .B1 (n_354), .B2 (n_353));
AND2_X1 i_415 (.ZN (n_351), .A1 (p_0[7]), .A2 (accumulator[7]));
NAND2_X1 i_414 (.ZN (n_350), .A1 (p_0[6]), .A2 (accumulator[6]));
INV_X1 i_413 (.ZN (n_349), .A (n_350));
NOR2_X1 i_412 (.ZN (n_348), .A1 (n_360), .A2 (n_350));
NOR4_X1 i_411 (.ZN (n_347), .A1 (n_351), .A2 (n_348), .A3 (n_352), .A4 (n_355));
NOR2_X1 i_410 (.ZN (n_346), .A1 (p_0[11]), .A2 (accumulator[11]));
NOR2_X1 i_409 (.ZN (n_345), .A1 (p_0[9]), .A2 (accumulator[9]));
NOR2_X1 i_408 (.ZN (n_344), .A1 (p_0[10]), .A2 (accumulator[10]));
OR3_X1 i_407 (.ZN (n_343), .A1 (n_346), .A2 (n_344), .A3 (n_345));
NOR2_X1 i_406 (.ZN (n_342), .A1 (p_0[8]), .A2 (accumulator[8]));
NOR3_X1 i_405 (.ZN (n_341), .A1 (n_343), .A2 (n_342), .A3 (n_347));
NAND2_X1 i_404 (.ZN (n_340), .A1 (p_0[8]), .A2 (accumulator[8]));
NAND2_X1 i_403 (.ZN (n_339), .A1 (p_0[9]), .A2 (accumulator[9]));
AOI21_X1 i_402 (.ZN (n_338), .A (n_343), .B1 (n_340), .B2 (n_339));
AND2_X1 i_401 (.ZN (n_337), .A1 (p_0[11]), .A2 (accumulator[11]));
NAND2_X1 i_400 (.ZN (n_336), .A1 (p_0[10]), .A2 (accumulator[10]));
INV_X1 i_399 (.ZN (n_335), .A (n_336));
NOR2_X1 i_398 (.ZN (n_334), .A1 (n_346), .A2 (n_336));
NOR4_X1 i_397 (.ZN (n_333), .A1 (n_337), .A2 (n_334), .A3 (n_338), .A4 (n_341));
NOR2_X1 i_396 (.ZN (n_332), .A1 (p_0[15]), .A2 (accumulator[15]));
NOR2_X1 i_395 (.ZN (n_331), .A1 (p_0[13]), .A2 (accumulator[13]));
NOR2_X1 i_394 (.ZN (n_330), .A1 (p_0[14]), .A2 (accumulator[14]));
OR3_X1 i_393 (.ZN (n_329), .A1 (n_332), .A2 (n_330), .A3 (n_331));
NOR2_X1 i_392 (.ZN (n_328), .A1 (p_0[12]), .A2 (accumulator[12]));
NOR3_X1 i_391 (.ZN (n_327), .A1 (n_329), .A2 (n_328), .A3 (n_333));
NAND2_X1 i_390 (.ZN (n_326), .A1 (p_0[12]), .A2 (accumulator[12]));
NAND2_X1 i_389 (.ZN (n_325), .A1 (p_0[13]), .A2 (accumulator[13]));
AOI21_X1 i_388 (.ZN (n_324), .A (n_329), .B1 (n_326), .B2 (n_325));
AND2_X1 i_387 (.ZN (n_323), .A1 (p_0[15]), .A2 (accumulator[15]));
NAND2_X1 i_386 (.ZN (n_322), .A1 (p_0[14]), .A2 (accumulator[14]));
INV_X1 i_385 (.ZN (n_321), .A (n_322));
NOR2_X1 i_384 (.ZN (n_320), .A1 (n_332), .A2 (n_322));
NOR4_X1 i_383 (.ZN (n_319), .A1 (n_323), .A2 (n_320), .A3 (n_324), .A4 (n_327));
NOR2_X1 i_382 (.ZN (n_318), .A1 (p_0[20]), .A2 (accumulator[20]));
NOR2_X1 i_381 (.ZN (n_317), .A1 (p_0[23]), .A2 (accumulator[23]));
INV_X1 i_380 (.ZN (n_316), .A (n_317));
NOR2_X1 i_379 (.ZN (n_315), .A1 (p_0[21]), .A2 (accumulator[21]));
INV_X1 i_378 (.ZN (n_314), .A (n_315));
NOR2_X1 i_377 (.ZN (n_313), .A1 (p_0[22]), .A2 (accumulator[22]));
INV_X1 i_376 (.ZN (n_312), .A (n_313));
NAND3_X1 i_375 (.ZN (n_311), .A1 (n_316), .A2 (n_312), .A3 (n_314));
OR2_X1 i_374 (.ZN (n_310), .A1 (n_318), .A2 (n_311));
NOR2_X1 i_373 (.ZN (n_309), .A1 (p_0[31]), .A2 (accumulator[31]));
INV_X1 i_372 (.ZN (n_308), .A (n_309));
NOR2_X1 i_371 (.ZN (n_307), .A1 (p_0[29]), .A2 (accumulator[29]));
INV_X1 i_370 (.ZN (n_306), .A (n_307));
NOR2_X1 i_369 (.ZN (n_305), .A1 (p_0[30]), .A2 (accumulator[30]));
INV_X1 i_368 (.ZN (n_304), .A (n_305));
NAND3_X1 i_367 (.ZN (n_303), .A1 (n_308), .A2 (n_304), .A3 (n_306));
NOR2_X1 i_366 (.ZN (n_302), .A1 (p_0[28]), .A2 (accumulator[28]));
OR2_X1 i_365 (.ZN (n_301), .A1 (n_303), .A2 (n_302));
NOR2_X1 i_364 (.ZN (n_300), .A1 (p_0[27]), .A2 (accumulator[27]));
INV_X1 i_363 (.ZN (n_299), .A (n_300));
NOR2_X1 i_362 (.ZN (n_298), .A1 (p_0[25]), .A2 (accumulator[25]));
INV_X1 i_361 (.ZN (n_297), .A (n_298));
NOR2_X1 i_360 (.ZN (n_296), .A1 (p_0[26]), .A2 (accumulator[26]));
INV_X1 i_359 (.ZN (n_295), .A (n_296));
NAND3_X1 i_358 (.ZN (n_294), .A1 (n_299), .A2 (n_295), .A3 (n_297));
NOR2_X1 i_357 (.ZN (n_293), .A1 (p_0[24]), .A2 (accumulator[24]));
OR2_X1 i_356 (.ZN (n_292), .A1 (n_294), .A2 (n_293));
OR2_X1 i_355 (.ZN (n_291), .A1 (n_301), .A2 (n_292));
OR2_X1 i_354 (.ZN (n_290), .A1 (n_310), .A2 (n_291));
NOR2_X1 i_353 (.ZN (n_289), .A1 (p_0[19]), .A2 (accumulator[19]));
INV_X1 i_352 (.ZN (n_288), .A (n_289));
NOR2_X1 i_351 (.ZN (n_287), .A1 (p_0[17]), .A2 (accumulator[17]));
INV_X1 i_350 (.ZN (n_286), .A (n_287));
NOR2_X1 i_349 (.ZN (n_285), .A1 (p_0[18]), .A2 (accumulator[18]));
INV_X1 i_348 (.ZN (n_284), .A (n_285));
NAND3_X1 i_347 (.ZN (n_283), .A1 (n_288), .A2 (n_284), .A3 (n_286));
NOR2_X1 i_346 (.ZN (n_282), .A1 (p_0[16]), .A2 (accumulator[16]));
OR2_X1 i_345 (.ZN (n_281), .A1 (n_283), .A2 (n_282));
NOR3_X1 i_344 (.ZN (n_280), .A1 (n_290), .A2 (n_281), .A3 (n_319));
NAND2_X1 i_343 (.ZN (n_279), .A1 (p_0[16]), .A2 (accumulator[16]));
NAND2_X1 i_342 (.ZN (n_278), .A1 (p_0[17]), .A2 (accumulator[17]));
INV_X1 i_341 (.ZN (n_277), .A (n_278));
AOI21_X1 i_340 (.ZN (n_276), .A (n_283), .B1 (n_279), .B2 (n_278));
AND2_X1 i_339 (.ZN (n_275), .A1 (p_0[18]), .A2 (accumulator[18]));
AOI221_X1 i_338 (.ZN (n_274), .A (n_276), .B1 (p_0[19]), .B2 (accumulator[19]), .C1 (n_288), .C2 (n_275));
NAND2_X1 i_337 (.ZN (n_273), .A1 (p_0[24]), .A2 (accumulator[24]));
NAND2_X1 i_336 (.ZN (n_272), .A1 (p_0[25]), .A2 (accumulator[25]));
INV_X1 i_335 (.ZN (n_271), .A (n_272));
AOI21_X1 i_334 (.ZN (n_270), .A (n_294), .B1 (n_273), .B2 (n_272));
AND2_X1 i_333 (.ZN (n_269), .A1 (p_0[26]), .A2 (accumulator[26]));
AOI221_X1 i_332 (.ZN (n_268), .A (n_270), .B1 (p_0[27]), .B2 (accumulator[27]), .C1 (n_299), .C2 (n_269));
NAND2_X1 i_331 (.ZN (n_267), .A1 (p_0[28]), .A2 (accumulator[28]));
AND2_X1 i_330 (.ZN (n_266), .A1 (p_0[29]), .A2 (accumulator[29]));
AOI21_X1 i_329 (.ZN (n_265), .A (n_266), .B1 (p_0[28]), .B2 (accumulator[28]));
NAND2_X1 i_328 (.ZN (n_264), .A1 (p_0[30]), .A2 (accumulator[30]));
INV_X1 i_327 (.ZN (n_263), .A (n_264));
OAI222_X1 i_326 (.ZN (n_262), .A1 (n_303), .A2 (n_265), .B1 (n_309), .B2 (n_264), .C1 (n_377), .C2 (n_373));
NAND2_X1 i_325 (.ZN (n_261), .A1 (p_0[20]), .A2 (accumulator[20]));
NAND2_X1 i_324 (.ZN (n_260), .A1 (p_0[21]), .A2 (accumulator[21]));
INV_X1 i_323 (.ZN (n_259), .A (n_260));
AOI21_X1 i_322 (.ZN (n_258), .A (n_311), .B1 (n_261), .B2 (n_260));
AND2_X1 i_321 (.ZN (n_257), .A1 (p_0[22]), .A2 (accumulator[22]));
AOI221_X1 i_320 (.ZN (n_256), .A (n_258), .B1 (p_0[23]), .B2 (accumulator[23]), .C1 (n_316), .C2 (n_257));
OAI222_X1 i_319 (.ZN (n_255), .A1 (n_290), .A2 (n_274), .B1 (n_291), .B2 (n_256), .C1 (n_301), .C2 (n_268));
NOR3_X1 i_318 (.ZN (n_254), .A1 (n_262), .A2 (n_255), .A3 (n_280));
NOR2_X1 i_317 (.ZN (n_253), .A1 (p_0[36]), .A2 (accumulator[36]));
NOR2_X1 i_316 (.ZN (n_252), .A1 (p_0[39]), .A2 (accumulator[39]));
INV_X1 i_315 (.ZN (n_251), .A (n_252));
NOR2_X1 i_314 (.ZN (n_250), .A1 (p_0[37]), .A2 (accumulator[37]));
INV_X1 i_313 (.ZN (n_249), .A (n_250));
NOR2_X1 i_312 (.ZN (n_248), .A1 (p_0[38]), .A2 (accumulator[38]));
INV_X1 i_311 (.ZN (n_247), .A (n_248));
NAND3_X1 i_310 (.ZN (n_246), .A1 (n_251), .A2 (n_247), .A3 (n_249));
OR2_X1 i_309 (.ZN (n_245), .A1 (n_253), .A2 (n_246));
NOR2_X1 i_308 (.ZN (n_244), .A1 (p_0[47]), .A2 (accumulator[47]));
NOR2_X1 i_307 (.ZN (n_243), .A1 (p_0[45]), .A2 (accumulator[45]));
NOR2_X1 i_306 (.ZN (n_242), .A1 (p_0[46]), .A2 (accumulator[46]));
NOR2_X1 i_305 (.ZN (n_241), .A1 (n_243), .A2 (n_242));
NOR3_X1 i_304 (.ZN (n_240), .A1 (n_244), .A2 (n_242), .A3 (n_243));
OAI21_X1 i_303 (.ZN (n_239), .A (n_240), .B1 (p_0[44]), .B2 (accumulator[44]));
NOR2_X1 i_302 (.ZN (n_238), .A1 (p_0[43]), .A2 (accumulator[43]));
INV_X1 i_301 (.ZN (n_237), .A (n_238));
NOR2_X1 i_300 (.ZN (n_236), .A1 (p_0[41]), .A2 (accumulator[41]));
INV_X1 i_299 (.ZN (n_235), .A (n_236));
NOR2_X1 i_298 (.ZN (n_234), .A1 (p_0[42]), .A2 (accumulator[42]));
INV_X1 i_297 (.ZN (n_233), .A (n_234));
NAND3_X1 i_296 (.ZN (n_232), .A1 (n_237), .A2 (n_233), .A3 (n_235));
NOR2_X1 i_295 (.ZN (n_231), .A1 (p_0[40]), .A2 (accumulator[40]));
OR2_X1 i_294 (.ZN (n_230), .A1 (n_232), .A2 (n_231));
OR2_X1 i_293 (.ZN (n_229), .A1 (n_239), .A2 (n_230));
OR2_X1 i_292 (.ZN (n_228), .A1 (n_245), .A2 (n_229));
NOR2_X1 i_291 (.ZN (n_227), .A1 (p_0[35]), .A2 (accumulator[35]));
INV_X1 i_290 (.ZN (n_226), .A (n_227));
NOR2_X1 i_289 (.ZN (n_225), .A1 (p_0[33]), .A2 (accumulator[33]));
INV_X1 i_288 (.ZN (n_224), .A (n_225));
NOR2_X1 i_287 (.ZN (n_223), .A1 (p_0[34]), .A2 (accumulator[34]));
INV_X1 i_286 (.ZN (n_222), .A (n_223));
NAND3_X1 i_285 (.ZN (n_221), .A1 (n_226), .A2 (n_222), .A3 (n_224));
NOR2_X1 i_284 (.ZN (n_220), .A1 (p_0[32]), .A2 (accumulator[32]));
OR2_X1 i_283 (.ZN (n_219), .A1 (n_221), .A2 (n_220));
NOR3_X1 i_282 (.ZN (n_218), .A1 (n_228), .A2 (n_219), .A3 (n_254));
NAND2_X1 i_281 (.ZN (n_217), .A1 (p_0[32]), .A2 (accumulator[32]));
NAND2_X1 i_280 (.ZN (n_216), .A1 (p_0[33]), .A2 (accumulator[33]));
INV_X1 i_279 (.ZN (n_215), .A (n_216));
AOI21_X1 i_278 (.ZN (n_214), .A (n_221), .B1 (n_217), .B2 (n_216));
AND2_X1 i_277 (.ZN (n_213), .A1 (p_0[34]), .A2 (accumulator[34]));
AOI221_X1 i_276 (.ZN (n_212), .A (n_214), .B1 (p_0[35]), .B2 (accumulator[35]), .C1 (n_226), .C2 (n_213));
NOR2_X1 i_275 (.ZN (n_211), .A1 (n_228), .A2 (n_212));
NAND2_X1 i_274 (.ZN (n_210), .A1 (p_0[36]), .A2 (accumulator[36]));
NAND2_X1 i_273 (.ZN (n_209), .A1 (p_0[37]), .A2 (accumulator[37]));
INV_X1 i_272 (.ZN (n_208), .A (n_209));
AOI21_X1 i_271 (.ZN (n_207), .A (n_246), .B1 (n_210), .B2 (n_209));
AND2_X1 i_270 (.ZN (n_206), .A1 (p_0[38]), .A2 (accumulator[38]));
AOI221_X1 i_269 (.ZN (n_205), .A (n_207), .B1 (p_0[39]), .B2 (accumulator[39]), .C1 (n_251), .C2 (n_206));
NAND2_X1 i_268 (.ZN (n_204), .A1 (p_0[44]), .A2 (accumulator[44]));
INV_X1 i_267 (.ZN (n_203), .A (n_204));
AND2_X1 i_266 (.ZN (n_202), .A1 (p_0[45]), .A2 (accumulator[45]));
OAI21_X1 i_265 (.ZN (n_201), .A (n_240), .B1 (n_203), .B2 (n_202));
NAND2_X1 i_264 (.ZN (n_200), .A1 (p_0[46]), .A2 (accumulator[46]));
INV_X1 i_263 (.ZN (n_199), .A (n_200));
OAI21_X1 i_262 (.ZN (n_198), .A (n_201), .B1 (n_244), .B2 (n_200));
AOI21_X1 i_261 (.ZN (n_197), .A (n_198), .B1 (p_0[47]), .B2 (accumulator[47]));
NAND2_X1 i_260 (.ZN (n_196), .A1 (p_0[40]), .A2 (accumulator[40]));
NAND2_X1 i_259 (.ZN (n_195), .A1 (p_0[41]), .A2 (accumulator[41]));
INV_X1 i_258 (.ZN (n_194), .A (n_195));
AOI21_X1 i_257 (.ZN (n_193), .A (n_232), .B1 (n_196), .B2 (n_195));
AND2_X1 i_256 (.ZN (n_192), .A1 (p_0[42]), .A2 (accumulator[42]));
AOI221_X1 i_255 (.ZN (n_191), .A (n_193), .B1 (p_0[43]), .B2 (accumulator[43]), .C1 (n_237), .C2 (n_192));
OAI221_X1 i_254 (.ZN (n_190), .A (n_197), .B1 (n_239), .B2 (n_191), .C1 (n_229), .C2 (n_205));
NOR3_X1 i_253 (.ZN (n_189), .A1 (n_211), .A2 (n_190), .A3 (n_218));
NOR2_X1 i_252 (.ZN (n_188), .A1 (p_0[51]), .A2 (accumulator[51]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (p_0[49]), .A2 (accumulator[49]));
NOR2_X1 i_250 (.ZN (n_186), .A1 (p_0[50]), .A2 (accumulator[50]));
OR3_X1 i_249 (.ZN (n_185), .A1 (n_188), .A2 (n_186), .A3 (n_187));
NOR2_X1 i_248 (.ZN (n_184), .A1 (p_0[48]), .A2 (accumulator[48]));
NOR3_X1 i_247 (.ZN (n_183), .A1 (n_185), .A2 (n_184), .A3 (n_189));
NAND2_X1 i_246 (.ZN (n_182), .A1 (p_0[48]), .A2 (accumulator[48]));
NAND2_X1 i_245 (.ZN (n_181), .A1 (p_0[49]), .A2 (accumulator[49]));
AOI21_X1 i_244 (.ZN (n_180), .A (n_185), .B1 (n_182), .B2 (n_181));
AND2_X1 i_243 (.ZN (n_179), .A1 (p_0[51]), .A2 (accumulator[51]));
NAND2_X1 i_242 (.ZN (n_178), .A1 (p_0[50]), .A2 (accumulator[50]));
INV_X1 i_241 (.ZN (n_177), .A (n_178));
NOR2_X1 i_240 (.ZN (n_176), .A1 (n_188), .A2 (n_178));
NOR4_X1 i_239 (.ZN (n_175), .A1 (n_179), .A2 (n_176), .A3 (n_180), .A4 (n_183));
NOR2_X1 i_238 (.ZN (n_174), .A1 (p_0[59]), .A2 (accumulator[59]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (p_0[57]), .A2 (accumulator[57]));
NOR2_X1 i_236 (.ZN (n_172), .A1 (p_0[58]), .A2 (accumulator[58]));
NOR2_X1 i_235 (.ZN (n_171), .A1 (n_173), .A2 (n_172));
NOR3_X1 i_234 (.ZN (n_170), .A1 (n_174), .A2 (n_172), .A3 (n_173));
OAI21_X1 i_233 (.ZN (n_169), .A (n_170), .B1 (p_0[56]), .B2 (accumulator[56]));
NOR2_X1 i_232 (.ZN (n_168), .A1 (p_0[55]), .A2 (accumulator[55]));
INV_X1 i_231 (.ZN (n_167), .A (n_168));
NOR2_X1 i_230 (.ZN (n_166), .A1 (p_0[53]), .A2 (accumulator[53]));
INV_X1 i_229 (.ZN (n_165), .A (n_166));
NOR2_X1 i_228 (.ZN (n_164), .A1 (p_0[54]), .A2 (accumulator[54]));
INV_X1 i_227 (.ZN (n_163), .A (n_164));
NAND3_X1 i_226 (.ZN (n_162), .A1 (n_167), .A2 (n_163), .A3 (n_165));
NOR2_X1 i_225 (.ZN (n_161), .A1 (p_0[52]), .A2 (accumulator[52]));
OR2_X1 i_224 (.ZN (n_160), .A1 (n_162), .A2 (n_161));
NOR3_X1 i_223 (.ZN (n_159), .A1 (n_169), .A2 (n_160), .A3 (n_175));
NAND2_X1 i_222 (.ZN (n_158), .A1 (p_0[52]), .A2 (accumulator[52]));
NAND2_X1 i_221 (.ZN (n_157), .A1 (p_0[53]), .A2 (accumulator[53]));
INV_X1 i_220 (.ZN (n_156), .A (n_157));
AOI21_X1 i_219 (.ZN (n_155), .A (n_162), .B1 (n_158), .B2 (n_157));
AND2_X1 i_218 (.ZN (n_154), .A1 (p_0[54]), .A2 (accumulator[54]));
AOI221_X1 i_217 (.ZN (n_153), .A (n_155), .B1 (p_0[55]), .B2 (accumulator[55]), .C1 (n_167), .C2 (n_154));
NOR2_X1 i_216 (.ZN (n_152), .A1 (n_169), .A2 (n_153));
NAND2_X1 i_215 (.ZN (n_151), .A1 (p_0[56]), .A2 (accumulator[56]));
INV_X1 i_214 (.ZN (n_150), .A (n_151));
AND2_X1 i_213 (.ZN (n_149), .A1 (p_0[57]), .A2 (accumulator[57]));
OAI21_X1 i_212 (.ZN (n_148), .A (n_170), .B1 (n_150), .B2 (n_149));
INV_X1 i_211 (.ZN (n_147), .A (n_148));
NAND2_X1 i_210 (.ZN (n_146), .A1 (p_0[58]), .A2 (accumulator[58]));
INV_X1 i_209 (.ZN (n_145), .A (n_146));
OAI22_X1 i_208 (.ZN (n_144), .A1 (n_378), .A2 (n_374), .B1 (n_174), .B2 (n_146));
NOR4_X1 i_207 (.ZN (n_143), .A1 (n_147), .A2 (n_144), .A3 (n_152), .A4 (n_159));
AOI21_X1 i_206 (.ZN (n_142), .A (n_371), .B1 (p_0[60]), .B2 (accumulator[60]));
AOI21_X1 i_205 (.ZN (n_141), .A (n_371), .B1 (n_143), .B2 (n_142));
INV_X1 i_204 (.ZN (n_140), .A (n_141));
NAND2_X1 i_203 (.ZN (n_139), .A1 (p_0[62]), .A2 (accumulator[62]));
INV_X1 i_202 (.ZN (n_138), .A (n_139));
NAND2_X1 i_201 (.ZN (n_137), .A1 (n_379), .A2 (n_375));
OAI21_X1 i_200 (.ZN (n_136), .A (n_137), .B1 (n_379), .B2 (n_375));
INV_X1 i_199 (.ZN (n_135), .A (n_136));
NAND3_X1 i_198 (.ZN (n_134), .A1 (n_139), .A2 (n_135), .A3 (n_140));
OAI221_X1 i_197 (.ZN (n_133), .A (n_134), .B1 (p_0[62]), .B2 (accumulator[62]), .C1 (n_138), .C2 (n_137));
XNOR2_X1 i_196 (.ZN (n_132), .A (p_0[63]), .B (accumulator[63]));
XOR2_X1 i_195 (.Z (p_1[63]), .A (n_133), .B (n_132));
OAI21_X1 i_194 (.ZN (n_131), .A (n_139), .B1 (p_0[62]), .B2 (accumulator[62]));
AOI22_X1 i_193 (.ZN (n_130), .A1 (p_0[61]), .A2 (accumulator[61]), .B1 (n_141), .B2 (n_137));
XOR2_X1 i_192 (.Z (p_1[62]), .A (n_131), .B (n_130));
AOI22_X1 i_191 (.ZN (p_1[61]), .A1 (n_140), .A2 (n_136), .B1 (n_141), .B2 (n_135));
XNOR2_X1 i_190 (.ZN (p_1[60]), .A (n_143), .B (n_142));
AOI21_X1 i_189 (.ZN (n_129), .A (n_174), .B1 (p_0[59]), .B2 (accumulator[59]));
OAI21_X1 i_188 (.ZN (n_128), .A (n_153), .B1 (n_175), .B2 (n_160));
OAI21_X1 i_187 (.ZN (n_127), .A (n_151), .B1 (p_0[56]), .B2 (accumulator[56]));
OAI22_X1 i_186 (.ZN (n_126), .A1 (p_0[56]), .A2 (accumulator[56]), .B1 (n_150), .B2 (n_128));
INV_X1 i_185 (.ZN (n_125), .A (n_126));
NOR2_X1 i_184 (.ZN (n_124), .A1 (n_173), .A2 (n_149));
NAND3_X1 i_183 (.ZN (n_123), .A1 (n_146), .A2 (n_124), .A3 (n_126));
OAI21_X1 i_182 (.ZN (n_122), .A (n_123), .B1 (n_171), .B2 (n_145));
XNOR2_X1 i_181 (.ZN (p_1[59]), .A (n_129), .B (n_122));
NOR2_X1 i_180 (.ZN (n_121), .A1 (n_172), .A2 (n_145));
OAI22_X1 i_179 (.ZN (n_120), .A1 (p_0[57]), .A2 (accumulator[57]), .B1 (n_149), .B2 (n_125));
XNOR2_X1 i_178 (.ZN (p_1[58]), .A (n_121), .B (n_120));
XOR2_X1 i_177 (.Z (p_1[57]), .A (n_125), .B (n_124));
XNOR2_X1 i_176 (.ZN (p_1[56]), .A (n_128), .B (n_127));
AOI21_X1 i_175 (.ZN (n_119), .A (n_168), .B1 (p_0[55]), .B2 (accumulator[55]));
OAI21_X1 i_174 (.ZN (n_118), .A (n_158), .B1 (p_0[52]), .B2 (accumulator[52]));
AOI21_X1 i_173 (.ZN (n_117), .A (n_161), .B1 (n_175), .B2 (n_158));
OAI21_X1 i_172 (.ZN (n_116), .A (n_165), .B1 (n_156), .B2 (n_117));
INV_X1 i_171 (.ZN (n_115), .A (n_116));
NOR2_X1 i_170 (.ZN (n_114), .A1 (n_166), .A2 (n_156));
OAI21_X1 i_169 (.ZN (n_113), .A (n_163), .B1 (n_154), .B2 (n_115));
XNOR2_X1 i_168 (.ZN (p_1[55]), .A (n_119), .B (n_113));
NOR2_X1 i_167 (.ZN (n_112), .A1 (n_164), .A2 (n_154));
XOR2_X1 i_166 (.Z (p_1[54]), .A (n_115), .B (n_112));
XOR2_X1 i_165 (.Z (p_1[53]), .A (n_117), .B (n_114));
XOR2_X1 i_164 (.Z (p_1[52]), .A (n_175), .B (n_118));
NOR2_X1 i_163 (.ZN (n_111), .A1 (n_188), .A2 (n_179));
OAI21_X1 i_162 (.ZN (n_110), .A (n_182), .B1 (p_0[48]), .B2 (accumulator[48]));
AOI21_X1 i_161 (.ZN (n_109), .A (n_184), .B1 (n_189), .B2 (n_182));
INV_X1 i_160 (.ZN (n_108), .A (n_109));
AOI21_X1 i_159 (.ZN (n_107), .A (n_187), .B1 (n_181), .B2 (n_108));
AOI21_X1 i_158 (.ZN (n_106), .A (n_187), .B1 (p_0[49]), .B2 (accumulator[49]));
OAI22_X1 i_157 (.ZN (n_105), .A1 (p_0[50]), .A2 (accumulator[50]), .B1 (n_177), .B2 (n_107));
XNOR2_X1 i_156 (.ZN (p_1[51]), .A (n_111), .B (n_105));
NOR2_X1 i_155 (.ZN (n_104), .A1 (n_186), .A2 (n_177));
XOR2_X1 i_154 (.Z (p_1[50]), .A (n_107), .B (n_104));
XOR2_X1 i_153 (.Z (p_1[49]), .A (n_109), .B (n_106));
XOR2_X1 i_152 (.Z (p_1[48]), .A (n_189), .B (n_110));
AOI21_X1 i_151 (.ZN (n_103), .A (n_244), .B1 (p_0[47]), .B2 (accumulator[47]));
OAI21_X1 i_150 (.ZN (n_102), .A (n_212), .B1 (n_254), .B2 (n_219));
INV_X1 i_149 (.ZN (n_101), .A (n_102));
OAI21_X1 i_148 (.ZN (n_100), .A (n_205), .B1 (n_245), .B2 (n_101));
INV_X1 i_147 (.ZN (n_99), .A (n_100));
OAI21_X1 i_146 (.ZN (n_98), .A (n_191), .B1 (n_230), .B2 (n_99));
OAI21_X1 i_145 (.ZN (n_97), .A (n_204), .B1 (p_0[44]), .B2 (accumulator[44]));
OAI22_X1 i_144 (.ZN (n_96), .A1 (p_0[44]), .A2 (accumulator[44]), .B1 (n_203), .B2 (n_98));
INV_X1 i_143 (.ZN (n_95), .A (n_96));
NOR2_X1 i_142 (.ZN (n_94), .A1 (n_243), .A2 (n_202));
NAND3_X1 i_141 (.ZN (n_93), .A1 (n_200), .A2 (n_94), .A3 (n_96));
OAI21_X1 i_140 (.ZN (n_92), .A (n_93), .B1 (n_241), .B2 (n_199));
XNOR2_X1 i_139 (.ZN (p_1[47]), .A (n_103), .B (n_92));
NOR2_X1 i_138 (.ZN (n_91), .A1 (n_242), .A2 (n_199));
OAI22_X1 i_137 (.ZN (n_90), .A1 (p_0[45]), .A2 (accumulator[45]), .B1 (n_202), .B2 (n_95));
XNOR2_X1 i_136 (.ZN (p_1[46]), .A (n_91), .B (n_90));
XOR2_X1 i_135 (.Z (p_1[45]), .A (n_95), .B (n_94));
XNOR2_X1 i_134 (.ZN (p_1[44]), .A (n_98), .B (n_97));
AOI21_X1 i_133 (.ZN (n_89), .A (n_238), .B1 (p_0[43]), .B2 (accumulator[43]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_196), .B1 (p_0[40]), .B2 (accumulator[40]));
AOI21_X1 i_131 (.ZN (n_87), .A (n_231), .B1 (n_196), .B2 (n_99));
OAI21_X1 i_130 (.ZN (n_86), .A (n_235), .B1 (n_194), .B2 (n_87));
INV_X1 i_129 (.ZN (n_85), .A (n_86));
NOR2_X1 i_128 (.ZN (n_84), .A1 (n_236), .A2 (n_194));
OAI21_X1 i_127 (.ZN (n_83), .A (n_233), .B1 (n_192), .B2 (n_85));
XNOR2_X1 i_126 (.ZN (p_1[43]), .A (n_89), .B (n_83));
NOR2_X1 i_125 (.ZN (n_82), .A1 (n_234), .A2 (n_192));
XOR2_X1 i_124 (.Z (p_1[42]), .A (n_85), .B (n_82));
XOR2_X1 i_123 (.Z (p_1[41]), .A (n_87), .B (n_84));
XOR2_X1 i_122 (.Z (p_1[40]), .A (n_99), .B (n_88));
AOI21_X1 i_121 (.ZN (n_81), .A (n_252), .B1 (p_0[39]), .B2 (accumulator[39]));
OAI21_X1 i_120 (.ZN (n_80), .A (n_210), .B1 (p_0[36]), .B2 (accumulator[36]));
AOI21_X1 i_119 (.ZN (n_79), .A (n_253), .B1 (n_210), .B2 (n_101));
OAI21_X1 i_118 (.ZN (n_78), .A (n_249), .B1 (n_208), .B2 (n_79));
INV_X1 i_117 (.ZN (n_77), .A (n_78));
NOR2_X1 i_116 (.ZN (n_76), .A1 (n_250), .A2 (n_208));
OAI21_X1 i_115 (.ZN (n_75), .A (n_247), .B1 (n_206), .B2 (n_77));
XNOR2_X1 i_114 (.ZN (p_1[39]), .A (n_81), .B (n_75));
NOR2_X1 i_113 (.ZN (n_74), .A1 (n_248), .A2 (n_206));
XOR2_X1 i_112 (.Z (p_1[38]), .A (n_77), .B (n_74));
XOR2_X1 i_111 (.Z (p_1[37]), .A (n_79), .B (n_76));
XOR2_X1 i_110 (.Z (p_1[36]), .A (n_101), .B (n_80));
AOI21_X1 i_109 (.ZN (n_73), .A (n_227), .B1 (p_0[35]), .B2 (accumulator[35]));
OAI21_X1 i_108 (.ZN (n_72), .A (n_217), .B1 (p_0[32]), .B2 (accumulator[32]));
AOI21_X1 i_107 (.ZN (n_71), .A (n_220), .B1 (n_254), .B2 (n_217));
OAI21_X1 i_106 (.ZN (n_70), .A (n_224), .B1 (n_215), .B2 (n_71));
INV_X1 i_105 (.ZN (n_69), .A (n_70));
NOR2_X1 i_104 (.ZN (n_68), .A1 (n_225), .A2 (n_215));
OAI21_X1 i_103 (.ZN (n_67), .A (n_222), .B1 (n_213), .B2 (n_69));
XNOR2_X1 i_102 (.ZN (p_1[35]), .A (n_73), .B (n_67));
NOR2_X1 i_101 (.ZN (n_66), .A1 (n_223), .A2 (n_213));
XOR2_X1 i_100 (.Z (p_1[34]), .A (n_69), .B (n_66));
XOR2_X1 i_99 (.Z (p_1[33]), .A (n_71), .B (n_68));
XOR2_X1 i_98 (.Z (p_1[32]), .A (n_254), .B (n_72));
OAI21_X1 i_97 (.ZN (n_65), .A (n_308), .B1 (n_377), .B2 (n_373));
OAI21_X1 i_96 (.ZN (n_64), .A (n_274), .B1 (n_319), .B2 (n_281));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
OAI21_X1 i_94 (.ZN (n_62), .A (n_256), .B1 (n_310), .B2 (n_63));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
OAI21_X1 i_92 (.ZN (n_60), .A (n_268), .B1 (n_292), .B2 (n_61));
INV_X1 i_91 (.ZN (n_59), .A (n_60));
OAI21_X1 i_90 (.ZN (n_58), .A (n_267), .B1 (p_0[28]), .B2 (accumulator[28]));
AOI21_X1 i_89 (.ZN (n_57), .A (n_302), .B1 (n_267), .B2 (n_59));
OAI21_X1 i_88 (.ZN (n_56), .A (n_306), .B1 (n_266), .B2 (n_57));
INV_X1 i_87 (.ZN (n_55), .A (n_56));
NOR2_X1 i_86 (.ZN (n_54), .A1 (n_307), .A2 (n_266));
OAI21_X1 i_85 (.ZN (n_53), .A (n_304), .B1 (n_263), .B2 (n_55));
XOR2_X1 i_84 (.Z (p_1[31]), .A (n_65), .B (n_53));
NOR2_X1 i_83 (.ZN (n_52), .A1 (n_305), .A2 (n_263));
XOR2_X1 i_82 (.Z (p_1[30]), .A (n_55), .B (n_52));
XOR2_X1 i_81 (.Z (p_1[29]), .A (n_57), .B (n_54));
XOR2_X1 i_80 (.Z (p_1[28]), .A (n_59), .B (n_58));
AOI21_X1 i_79 (.ZN (n_51), .A (n_300), .B1 (p_0[27]), .B2 (accumulator[27]));
OAI21_X1 i_78 (.ZN (n_50), .A (n_273), .B1 (p_0[24]), .B2 (accumulator[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_293), .B1 (n_273), .B2 (n_61));
OAI21_X1 i_76 (.ZN (n_48), .A (n_297), .B1 (n_271), .B2 (n_49));
INV_X1 i_75 (.ZN (n_47), .A (n_48));
NOR2_X1 i_74 (.ZN (n_46), .A1 (n_298), .A2 (n_271));
OAI21_X1 i_73 (.ZN (n_45), .A (n_295), .B1 (n_269), .B2 (n_47));
XNOR2_X1 i_72 (.ZN (p_1[27]), .A (n_51), .B (n_45));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_296), .A2 (n_269));
XOR2_X1 i_70 (.Z (p_1[26]), .A (n_47), .B (n_44));
XOR2_X1 i_69 (.Z (p_1[25]), .A (n_49), .B (n_46));
XOR2_X1 i_68 (.Z (p_1[24]), .A (n_61), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_317), .B1 (p_0[23]), .B2 (accumulator[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_261), .B1 (p_0[20]), .B2 (accumulator[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_318), .B1 (n_261), .B2 (n_63));
OAI21_X1 i_64 (.ZN (n_40), .A (n_314), .B1 (n_259), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_315), .A2 (n_259));
OAI21_X1 i_61 (.ZN (n_37), .A (n_312), .B1 (n_257), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_313), .A2 (n_257));
XOR2_X1 i_58 (.Z (p_1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_1[20]), .A (n_63), .B (n_42));
AOI21_X1 i_55 (.ZN (n_35), .A (n_289), .B1 (p_0[19]), .B2 (accumulator[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_279), .B1 (p_0[16]), .B2 (accumulator[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_282), .B1 (n_319), .B2 (n_279));
OAI21_X1 i_52 (.ZN (n_32), .A (n_286), .B1 (n_277), .B2 (n_33));
INV_X1 i_51 (.ZN (n_31), .A (n_32));
NOR2_X1 i_50 (.ZN (n_30), .A1 (n_287), .A2 (n_277));
OAI21_X1 i_49 (.ZN (n_29), .A (n_284), .B1 (n_275), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_285), .A2 (n_275));
XOR2_X1 i_46 (.Z (p_1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_1[16]), .A (n_319), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_332), .A2 (n_323));
OAI21_X1 i_42 (.ZN (n_26), .A (n_326), .B1 (p_0[12]), .B2 (accumulator[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_328), .B1 (n_333), .B2 (n_326));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_331), .B1 (n_325), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_331), .B1 (p_0[13]), .B2 (accumulator[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (accumulator[14]), .B1 (n_321), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_330), .A2 (n_321));
XOR2_X1 i_34 (.Z (p_1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_1[12]), .A (n_333), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_346), .A2 (n_337));
AOI21_X1 i_30 (.ZN (n_18), .A (n_342), .B1 (p_0[8]), .B2 (accumulator[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_342), .B1 (n_347), .B2 (n_340));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_345), .B1 (n_339), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_345), .B1 (p_0[9]), .B2 (accumulator[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (accumulator[10]), .B1 (n_335), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_344), .A2 (n_335));
XOR2_X1 i_22 (.Z (p_1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_1[8]), .A (n_347), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_360), .A2 (n_351));
OAI21_X1 i_18 (.ZN (n_10), .A (n_354), .B1 (p_0[4]), .B2 (accumulator[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_356), .B1 (n_361), .B2 (n_354));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_359), .B1 (n_353), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_359), .B1 (p_0[5]), .B2 (accumulator[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (accumulator[6]), .B1 (n_349), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_358), .A2 (n_349));
XOR2_X1 i_10 (.Z (p_1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_1[4]), .A (n_361), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_370), .B1 (n_376), .B2 (n_372));
XOR2_X1 i_6 (.Z (p_1[3]), .A (n_363), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_369), .B1 (p_0[2]), .B2 (accumulator[2]));
XNOR2_X1 i_4 (.ZN (p_1[2]), .A (n_364), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_365), .B1 (p_0[1]), .B2 (spw_n22));
XOR2_X1 i_2 (.Z (p_1[1]), .A (n_366), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_366), .B1 (p_0[0]), .B2 (spw_n8));
INV_X1 i_0 (.ZN (p_1[0]), .A (n_0));
CLKBUF_X1 spw__L2_c3_c1 (.Z (spw_n8), .A (accumulator[0]));
CLKBUF_X1 spw__L2_c2_c4 (.Z (spw_n22), .A (spw__n11));
CLKBUF_X1 spw__L2_c3_c5 (.Z (spw__n10), .A (spw__n11));
CLKBUF_X1 spw__L1_c1_c6 (.Z (spw__n11), .A (accumulator[1]));

endmodule //datapath__0_15

module datapath__0_12 (p_0, multiplicand_reg);

output [31:0] p_0;
input [31:0] multiplicand_reg;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (multiplicand_reg[25]));
INV_X1 i_63 (.ZN (n_32), .A (multiplicand_reg[21]));
INV_X1 i_62 (.ZN (n_31), .A (multiplicand_reg[14]));
INV_X1 i_61 (.ZN (n_30), .A (multiplicand_reg[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (multiplicand_reg[2]), .A2 (multiplicand_reg[1]), .A3 (multiplicand_reg[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (multiplicand_reg[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (multiplicand_reg[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (multiplicand_reg[5]), .A3 (multiplicand_reg[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (multiplicand_reg[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (multiplicand_reg[8]), .A3 (multiplicand_reg[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (multiplicand_reg[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (multiplicand_reg[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (multiplicand_reg[12]), .A3 (multiplicand_reg[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (multiplicand_reg[15]), .A3 (multiplicand_reg[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (multiplicand_reg[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (multiplicand_reg[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (multiplicand_reg[18]), .A3 (multiplicand_reg[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (multiplicand_reg[18]), .A3 (multiplicand_reg[19]), .A4 (multiplicand_reg[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (multiplicand_reg[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (multiplicand_reg[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (multiplicand_reg[23]), .A3 (multiplicand_reg[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (multiplicand_reg[26]), .A3 (multiplicand_reg[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (multiplicand_reg[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (multiplicand_reg[28]), .A3 (multiplicand_reg[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (multiplicand_reg[28]), .A3 (multiplicand_reg[29]), .A4 (multiplicand_reg[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (multiplicand_reg[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (multiplicand_reg[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (multiplicand_reg[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (multiplicand_reg[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (multiplicand_reg[27]), .B1 (n_9), .B2 (multiplicand_reg[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (multiplicand_reg[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (multiplicand_reg[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (multiplicand_reg[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (multiplicand_reg[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (multiplicand_reg[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (multiplicand_reg[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (multiplicand_reg[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (multiplicand_reg[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (multiplicand_reg[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (multiplicand_reg[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (multiplicand_reg[16]), .B1 (n_19), .B2 (multiplicand_reg[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (multiplicand_reg[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (multiplicand_reg[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (multiplicand_reg[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (multiplicand_reg[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (multiplicand_reg[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (multiplicand_reg[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (multiplicand_reg[9]), .B1 (n_25), .B2 (multiplicand_reg[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (multiplicand_reg[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (multiplicand_reg[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (multiplicand_reg[6]), .B1 (n_27), .B2 (multiplicand_reg[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (multiplicand_reg[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (multiplicand_reg[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (multiplicand_reg[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (multiplicand_reg[2]), .B1 (multiplicand_reg[1]), .B2 (multiplicand_reg[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (multiplicand_reg[1]), .B (multiplicand_reg[0]));

endmodule //datapath__0_12

module datapath__0_3 (p_0, multiplier_reg);

output [31:0] p_0;
input [31:0] multiplier_reg;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (multiplier_reg[25]));
INV_X1 i_63 (.ZN (n_32), .A (multiplier_reg[21]));
INV_X1 i_62 (.ZN (n_31), .A (multiplier_reg[14]));
INV_X1 i_61 (.ZN (n_30), .A (multiplier_reg[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (multiplier_reg[2]), .A2 (multiplier_reg[1]), .A3 (multiplier_reg[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (multiplier_reg[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (multiplier_reg[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (multiplier_reg[5]), .A3 (multiplier_reg[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (multiplier_reg[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (multiplier_reg[8]), .A3 (multiplier_reg[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (multiplier_reg[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (multiplier_reg[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (multiplier_reg[12]), .A3 (multiplier_reg[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (multiplier_reg[15]), .A3 (multiplier_reg[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (multiplier_reg[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (multiplier_reg[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (multiplier_reg[18]), .A3 (multiplier_reg[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (multiplier_reg[18]), .A3 (multiplier_reg[19]), .A4 (multiplier_reg[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (multiplier_reg[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (multiplier_reg[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (multiplier_reg[23]), .A3 (multiplier_reg[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (multiplier_reg[26]), .A3 (multiplier_reg[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (multiplier_reg[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (multiplier_reg[28]), .A3 (multiplier_reg[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (multiplier_reg[28]), .A3 (multiplier_reg[29]), .A4 (multiplier_reg[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (multiplier_reg[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (multiplier_reg[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (multiplier_reg[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (multiplier_reg[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (multiplier_reg[27]), .B1 (n_9), .B2 (multiplier_reg[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (multiplier_reg[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (multiplier_reg[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (multiplier_reg[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (multiplier_reg[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (multiplier_reg[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (multiplier_reg[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (multiplier_reg[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (multiplier_reg[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (multiplier_reg[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (multiplier_reg[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (multiplier_reg[16]), .B1 (n_19), .B2 (multiplier_reg[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (multiplier_reg[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (multiplier_reg[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (multiplier_reg[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (multiplier_reg[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (multiplier_reg[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (multiplier_reg[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (multiplier_reg[9]), .B1 (n_25), .B2 (multiplier_reg[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (multiplier_reg[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (multiplier_reg[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (multiplier_reg[6]), .B1 (n_27), .B2 (multiplier_reg[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (multiplier_reg[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (multiplier_reg[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (multiplier_reg[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (multiplier_reg[2]), .B1 (multiplier_reg[1]), .B2 (multiplier_reg[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (multiplier_reg[1]), .B (multiplier_reg[0]));

endmodule //datapath__0_3

module datapath (accumulator_0_PP_0, accumulator_1_PP_0, p_0, accumulator);

output [63:0] p_0;
input [63:0] accumulator;
input accumulator_0_PP_0;
input accumulator_1_PP_0;
wire spw_n156;
wire n_61;
wire n_0;
wire n_60;
wire n_59;
wire n_58;
wire n_1;
wire n_57;
wire n_56;
wire n_2;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_3;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_4;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_5;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire spt__n1;
wire spw__n227;


INV_X1 i_135 (.ZN (n_72), .A (accumulator[60]));
INV_X1 i_134 (.ZN (n_71), .A (accumulator[55]));
INV_X1 i_133 (.ZN (n_70), .A (accumulator[51]));
INV_X1 i_132 (.ZN (n_69), .A (accumulator[42]));
INV_X1 i_131 (.ZN (n_68), .A (accumulator[40]));
INV_X1 i_130 (.ZN (n_67), .A (accumulator[36]));
INV_X1 i_129 (.ZN (n_66), .A (accumulator[31]));
INV_X1 i_128 (.ZN (n_65), .A (accumulator[26]));
INV_X1 i_127 (.ZN (n_64), .A (accumulator[21]));
INV_X1 i_126 (.ZN (n_63), .A (accumulator[13]));
INV_X1 i_125 (.ZN (n_62), .A (accumulator[11]));
OR3_X4 i_124 (.ZN (n_61), .A1 (accumulator[2]), .A2 (accumulator[1]), .A3 (accumulator_0_PP_0));
OR2_X4 i_123 (.ZN (n_60), .A1 (n_61), .A2 (accumulator[3]));
OR2_X4 i_122 (.ZN (n_59), .A1 (n_60), .A2 (accumulator[4]));
OR3_X4 i_121 (.ZN (n_58), .A1 (n_59), .A2 (accumulator[5]), .A3 (accumulator[6]));
OR2_X4 i_120 (.ZN (n_57), .A1 (n_58), .A2 (accumulator[7]));
OR3_X4 i_119 (.ZN (n_56), .A1 (n_57), .A2 (accumulator[8]), .A3 (accumulator[9]));
NOR2_X4 i_118 (.ZN (n_55), .A1 (n_56), .A2 (accumulator[10]));
NAND2_X4 i_117 (.ZN (n_54), .A1 (n_55), .A2 (n_62));
NOR2_X4 i_116 (.ZN (n_53), .A1 (n_54), .A2 (accumulator[12]));
NAND2_X4 i_115 (.ZN (n_52), .A1 (n_53), .A2 (n_63));
OR3_X4 i_114 (.ZN (n_51), .A1 (n_52), .A2 (accumulator[14]), .A3 (accumulator[15]));
OR2_X4 i_113 (.ZN (n_50), .A1 (n_51), .A2 (accumulator[16]));
OR2_X4 i_112 (.ZN (n_49), .A1 (n_50), .A2 (accumulator[17]));
NOR2_X1 i_111 (.ZN (n_48), .A1 (n_49), .A2 (accumulator[18]));
NOR3_X1 i_110 (.ZN (n_47), .A1 (n_49), .A2 (accumulator[18]), .A3 (accumulator[19]));
NOR4_X4 i_109 (.ZN (n_46), .A1 (n_49), .A2 (accumulator[18]), .A3 (accumulator[19]), .A4 (accumulator[20]));
NAND2_X2 i_108 (.ZN (n_45), .A1 (n_46), .A2 (n_64));
OR2_X4 i_107 (.ZN (n_44), .A1 (n_45), .A2 (accumulator[22]));
NOR2_X1 i_106 (.ZN (n_43), .A1 (n_44), .A2 (accumulator[23]));
NOR3_X1 i_105 (.ZN (n_42), .A1 (n_44), .A2 (accumulator[23]), .A3 (accumulator[24]));
NOR4_X4 i_104 (.ZN (n_41), .A1 (n_44), .A2 (accumulator[23]), .A3 (accumulator[24]), .A4 (accumulator[25]));
NAND2_X2 i_103 (.ZN (n_40), .A1 (n_41), .A2 (n_65));
OR2_X4 i_102 (.ZN (n_39), .A1 (n_40), .A2 (accumulator[27]));
NOR2_X1 i_101 (.ZN (n_38), .A1 (n_39), .A2 (accumulator[28]));
NOR3_X1 i_100 (.ZN (n_37), .A1 (n_39), .A2 (accumulator[28]), .A3 (accumulator[29]));
NOR4_X4 i_99 (.ZN (n_36), .A1 (n_39), .A2 (accumulator[28]), .A3 (accumulator[29]), .A4 (accumulator[30]));
NAND2_X2 i_98 (.ZN (n_35), .A1 (n_36), .A2 (n_66));
OR2_X4 i_97 (.ZN (n_34), .A1 (n_35), .A2 (accumulator[32]));
NOR2_X1 i_96 (.ZN (n_33), .A1 (spw__n227), .A2 (accumulator[33]));
NOR3_X1 i_95 (.ZN (n_32), .A1 (spw__n227), .A2 (accumulator[33]), .A3 (accumulator[34]));
NOR4_X4 i_94 (.ZN (spt__n1), .A1 (n_34), .A2 (accumulator[33]), .A3 (accumulator[34]), .A4 (accumulator[35]));
NAND2_X2 i_93 (.ZN (n_30), .A1 (spt__n1), .A2 (n_67));
OR2_X4 i_92 (.ZN (n_29), .A1 (n_30), .A2 (accumulator[37]));
NOR2_X1 i_91 (.ZN (n_28), .A1 (n_29), .A2 (accumulator[38]));
NOR3_X4 i_90 (.ZN (n_27), .A1 (n_29), .A2 (accumulator[38]), .A3 (accumulator[39]));
NAND2_X2 i_89 (.ZN (n_26), .A1 (n_27), .A2 (n_68));
NOR2_X4 i_88 (.ZN (n_25), .A1 (n_26), .A2 (accumulator[41]));
NAND2_X2 i_87 (.ZN (n_24), .A1 (n_25), .A2 (n_69));
OR3_X4 i_86 (.ZN (n_23), .A1 (n_24), .A2 (accumulator[43]), .A3 (accumulator[44]));
OR2_X4 i_85 (.ZN (n_22), .A1 (n_23), .A2 (accumulator[45]));
OR2_X4 i_84 (.ZN (n_21), .A1 (n_22), .A2 (accumulator[46]));
OR2_X4 i_83 (.ZN (n_20), .A1 (n_21), .A2 (accumulator[47]));
NOR2_X1 i_82 (.ZN (n_19), .A1 (n_20), .A2 (accumulator[48]));
NOR3_X1 i_81 (.ZN (n_18), .A1 (n_20), .A2 (accumulator[48]), .A3 (accumulator[49]));
NOR4_X4 i_80 (.ZN (n_17), .A1 (n_20), .A2 (accumulator[48]), .A3 (accumulator[49]), .A4 (accumulator[50]));
NAND2_X4 i_79 (.ZN (n_16), .A1 (n_17), .A2 (n_70));
NOR2_X1 i_78 (.ZN (n_15), .A1 (n_16), .A2 (accumulator[52]));
NOR3_X1 i_77 (.ZN (n_14), .A1 (n_16), .A2 (accumulator[52]), .A3 (accumulator[53]));
NOR4_X4 i_76 (.ZN (n_13), .A1 (n_16), .A2 (accumulator[52]), .A3 (accumulator[53]), .A4 (accumulator[54]));
NAND2_X2 i_75 (.ZN (n_12), .A1 (n_13), .A2 (n_71));
OR3_X4 i_74 (.ZN (n_11), .A1 (n_12), .A2 (accumulator[56]), .A3 (accumulator[57]));
NOR2_X1 i_73 (.ZN (n_10), .A1 (n_11), .A2 (accumulator[58]));
NOR3_X4 i_72 (.ZN (n_9), .A1 (n_11), .A2 (accumulator[58]), .A3 (accumulator[59]));
NAND2_X4 i_71 (.ZN (n_8), .A1 (n_9), .A2 (n_72));
NOR2_X2 i_70 (.ZN (n_7), .A1 (n_8), .A2 (accumulator[61]));
NOR3_X4 i_69 (.ZN (n_6), .A1 (n_8), .A2 (accumulator[61]), .A3 (accumulator[62]));
XNOR2_X1 i_68 (.ZN (p_0[63]), .A (accumulator[63]), .B (n_6));
XNOR2_X1 i_67 (.ZN (p_0[62]), .A (accumulator[62]), .B (n_7));
XOR2_X1 i_66 (.Z (p_0[61]), .A (accumulator[61]), .B (n_8));
XNOR2_X1 i_65 (.ZN (p_0[60]), .A (accumulator[60]), .B (n_9));
XNOR2_X1 i_64 (.ZN (p_0[59]), .A (accumulator[59]), .B (n_10));
XOR2_X1 i_63 (.Z (p_0[58]), .A (accumulator[58]), .B (n_11));
OAI21_X1 i_62 (.ZN (n_5), .A (accumulator[57]), .B1 (n_12), .B2 (accumulator[56]));
AND2_X1 i_61 (.ZN (p_0[57]), .A1 (n_11), .A2 (n_5));
XOR2_X1 i_60 (.Z (p_0[56]), .A (accumulator[56]), .B (n_12));
XNOR2_X1 i_59 (.ZN (p_0[55]), .A (accumulator[55]), .B (n_13));
XNOR2_X1 i_58 (.ZN (p_0[54]), .A (accumulator[54]), .B (n_14));
XNOR2_X1 i_57 (.ZN (p_0[53]), .A (accumulator[53]), .B (n_15));
XOR2_X1 i_56 (.Z (p_0[52]), .A (accumulator[52]), .B (n_16));
XNOR2_X1 i_55 (.ZN (p_0[51]), .A (accumulator[51]), .B (n_17));
XNOR2_X1 i_54 (.ZN (p_0[50]), .A (accumulator[50]), .B (n_18));
XNOR2_X1 i_53 (.ZN (p_0[49]), .A (accumulator[49]), .B (n_19));
XOR2_X1 i_52 (.Z (p_0[48]), .A (accumulator[48]), .B (n_20));
XOR2_X1 i_51 (.Z (p_0[47]), .A (accumulator[47]), .B (n_21));
XOR2_X1 i_50 (.Z (p_0[46]), .A (accumulator[46]), .B (n_22));
XOR2_X1 i_49 (.Z (p_0[45]), .A (accumulator[45]), .B (n_23));
OAI21_X1 i_48 (.ZN (n_4), .A (accumulator[44]), .B1 (n_24), .B2 (accumulator[43]));
AND2_X1 i_47 (.ZN (p_0[44]), .A1 (n_23), .A2 (n_4));
XOR2_X1 i_46 (.Z (p_0[43]), .A (accumulator[43]), .B (n_24));
XNOR2_X1 i_45 (.ZN (p_0[42]), .A (accumulator[42]), .B (n_25));
XOR2_X1 i_44 (.Z (p_0[41]), .A (accumulator[41]), .B (n_26));
XNOR2_X1 i_43 (.ZN (p_0[40]), .A (accumulator[40]), .B (n_27));
XNOR2_X1 i_42 (.ZN (p_0[39]), .A (accumulator[39]), .B (n_28));
XOR2_X1 i_41 (.Z (p_0[38]), .A (accumulator[38]), .B (n_29));
XOR2_X1 i_40 (.Z (p_0[37]), .A (accumulator[37]), .B (n_30));
XNOR2_X1 i_39 (.ZN (p_0[36]), .A (accumulator[36]), .B (spt__n1));
XNOR2_X1 i_38 (.ZN (p_0[35]), .A (accumulator[35]), .B (n_32));
XNOR2_X1 i_37 (.ZN (p_0[34]), .A (accumulator[34]), .B (n_33));
XOR2_X1 i_36 (.Z (p_0[33]), .A (accumulator[33]), .B (n_34));
XOR2_X1 i_35 (.Z (p_0[32]), .A (accumulator[32]), .B (n_35));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (accumulator[31]), .B (n_36));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (accumulator[30]), .B (n_37));
XNOR2_X1 i_32 (.ZN (p_0[29]), .A (accumulator[29]), .B (n_38));
XOR2_X1 i_31 (.Z (p_0[28]), .A (accumulator[28]), .B (n_39));
XOR2_X1 i_30 (.Z (p_0[27]), .A (accumulator[27]), .B (n_40));
XNOR2_X1 i_29 (.ZN (p_0[26]), .A (accumulator[26]), .B (n_41));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (accumulator[25]), .B (n_42));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (accumulator[24]), .B (n_43));
XOR2_X1 i_26 (.Z (p_0[23]), .A (accumulator[23]), .B (n_44));
XOR2_X1 i_25 (.Z (p_0[22]), .A (accumulator[22]), .B (n_45));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (accumulator[21]), .B (n_46));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (accumulator[20]), .B (n_47));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (accumulator[19]), .B (n_48));
XOR2_X1 i_21 (.Z (p_0[18]), .A (accumulator[18]), .B (n_49));
XOR2_X1 i_20 (.Z (p_0[17]), .A (accumulator[17]), .B (n_50));
XOR2_X1 i_19 (.Z (p_0[16]), .A (accumulator[16]), .B (n_51));
OAI21_X1 i_18 (.ZN (n_3), .A (accumulator[15]), .B1 (n_52), .B2 (accumulator[14]));
AND2_X1 i_17 (.ZN (p_0[15]), .A1 (n_51), .A2 (n_3));
XOR2_X1 i_16 (.Z (p_0[14]), .A (accumulator[14]), .B (n_52));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (accumulator[13]), .B (n_53));
XOR2_X1 i_14 (.Z (p_0[12]), .A (accumulator[12]), .B (n_54));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (accumulator[11]), .B (n_55));
XOR2_X1 i_12 (.Z (p_0[10]), .A (accumulator[10]), .B (n_56));
OAI21_X1 i_11 (.ZN (n_2), .A (accumulator[9]), .B1 (n_57), .B2 (accumulator[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_56), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (accumulator[8]), .B (n_57));
XOR2_X1 i_8 (.Z (p_0[7]), .A (accumulator[7]), .B (n_58));
OAI21_X1 i_7 (.ZN (n_1), .A (accumulator[6]), .B1 (n_59), .B2 (accumulator[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_58), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (accumulator[5]), .B (n_59));
XOR2_X1 i_4 (.Z (p_0[4]), .A (accumulator[4]), .B (n_60));
XOR2_X1 i_3 (.Z (p_0[3]), .A (accumulator[3]), .B (n_61));
OAI21_X1 i_2 (.ZN (n_0), .A (accumulator[2]), .B1 (accumulator[1]), .B2 (accumulator_0_PP_0));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_61), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (spw_n156), .B (accumulator[0]));
CLKBUF_X1 spw__L1_c4_c125 (.Z (spw_n156), .A (accumulator_1_PP_0));
CLKBUF_X1 spw__L1_c197 (.Z (spw__n227), .A (n_34));

endmodule //datapath

module registerNbits (clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits

module registerNbits__0_28 (clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits__0_28

module registerNbits__0_25 (clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire spc__n1;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (spc__n1), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));
BUF_X8 spc__L1_c1_c1 (.Z (out[31]), .A (spc__n1));

endmodule //registerNbits__0_25

module registerNbits__0_22 (clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire spc__n1;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (spc__n1), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));
BUF_X8 spc__L1_c1_c1 (.Z (out[31]), .A (spc__n1));

endmodule //registerNbits__0_22

module sequential_multiplier (clk, set_signal, multipicand, multiplier, product, 
    reset, en);

output [63:0] product;
input clk;
input en;
input [31:0] multipicand;
input [31:0] multiplier;
input reset;
input set_signal;
wire \multiplicand_reg[31] ;
wire \multiplicand_reg[30] ;
wire \multiplicand_reg[29] ;
wire \multiplicand_reg[28] ;
wire \multiplicand_reg[27] ;
wire \multiplicand_reg[26] ;
wire \multiplicand_reg[25] ;
wire \multiplicand_reg[24] ;
wire \multiplicand_reg[23] ;
wire \multiplicand_reg[22] ;
wire \multiplicand_reg[21] ;
wire \multiplicand_reg[20] ;
wire \multiplicand_reg[19] ;
wire \multiplicand_reg[18] ;
wire \multiplicand_reg[17] ;
wire \multiplicand_reg[16] ;
wire \multiplicand_reg[15] ;
wire \multiplicand_reg[14] ;
wire \multiplicand_reg[13] ;
wire \multiplicand_reg[12] ;
wire \multiplicand_reg[11] ;
wire \multiplicand_reg[10] ;
wire \multiplicand_reg[9] ;
wire \multiplicand_reg[8] ;
wire \multiplicand_reg[7] ;
wire \multiplicand_reg[6] ;
wire \multiplicand_reg[5] ;
wire \multiplicand_reg[4] ;
wire \multiplicand_reg[3] ;
wire \multiplicand_reg[2] ;
wire \multiplicand_reg[1] ;
wire \multiplicand_reg[0] ;
wire \multiplier_reg[31] ;
wire \multiplier_reg[30] ;
wire \multiplier_reg[29] ;
wire \multiplier_reg[28] ;
wire \multiplier_reg[27] ;
wire \multiplier_reg[26] ;
wire \multiplier_reg[25] ;
wire \multiplier_reg[24] ;
wire \multiplier_reg[23] ;
wire \multiplier_reg[22] ;
wire \multiplier_reg[21] ;
wire \multiplier_reg[20] ;
wire \multiplier_reg[19] ;
wire \multiplier_reg[18] ;
wire \multiplier_reg[17] ;
wire \multiplier_reg[16] ;
wire \multiplier_reg[15] ;
wire \multiplier_reg[14] ;
wire \multiplier_reg[13] ;
wire \multiplier_reg[12] ;
wire \multiplier_reg[11] ;
wire \multiplier_reg[10] ;
wire \multiplier_reg[9] ;
wire \multiplier_reg[8] ;
wire \multiplier_reg[7] ;
wire \multiplier_reg[6] ;
wire \multiplier_reg[5] ;
wire \multiplier_reg[4] ;
wire \multiplier_reg[3] ;
wire \multiplier_reg[2] ;
wire \multiplier_reg[1] ;
wire \multiplier_reg[0] ;
wire \outmultiplier_reg[31] ;
wire \outmultiplier_reg[30] ;
wire \outmultiplier_reg[29] ;
wire \outmultiplier_reg[28] ;
wire \outmultiplier_reg[27] ;
wire \outmultiplier_reg[26] ;
wire \outmultiplier_reg[25] ;
wire \outmultiplier_reg[24] ;
wire \outmultiplier_reg[23] ;
wire \outmultiplier_reg[22] ;
wire \outmultiplier_reg[21] ;
wire \outmultiplier_reg[20] ;
wire \outmultiplier_reg[19] ;
wire \outmultiplier_reg[18] ;
wire \outmultiplier_reg[17] ;
wire \outmultiplier_reg[16] ;
wire \outmultiplier_reg[15] ;
wire \outmultiplier_reg[14] ;
wire \outmultiplier_reg[13] ;
wire \outmultiplier_reg[12] ;
wire \outmultiplier_reg[11] ;
wire \outmultiplier_reg[10] ;
wire \outmultiplier_reg[9] ;
wire \outmultiplier_reg[8] ;
wire \outmultiplier_reg[7] ;
wire \outmultiplier_reg[6] ;
wire \outmultiplier_reg[5] ;
wire \outmultiplier_reg[4] ;
wire \outmultiplier_reg[3] ;
wire \outmultiplier_reg[2] ;
wire \outmultiplier_reg[1] ;
wire \outmultiplier_reg[0] ;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_2_4;
wire n_0_2_0;
wire n_0_2_5;
wire n_0_2_1;
wire n_0_2_6;
wire n_0_2_2;
wire n_0_2_7;
wire n_0_2_3;
wire n_0_255;
wire n_0_2_8;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_2_9;
wire n_0_2_10;
wire n_0_324;
wire n_0_2_11;
wire n_0_2_12;
wire n_0_2_13;
wire n_0_2_14;
wire n_0_2_15;
wire n_0_453;
wire n_0_2_16;
wire n_0_2_17;
wire n_0_325;
wire n_0_2_18;
wire n_0_2_19;
wire n_0_390;
wire n_0_2_20;
wire n_0_2_21;
wire n_0_2_22;
wire n_0_326;
wire n_0_2_23;
wire n_0_391;
wire n_0_2_24;
wire n_0_327;
wire n_0_2_25;
wire n_0_392;
wire n_0_2_26;
wire n_0_328;
wire n_0_2_27;
wire n_0_393;
wire n_0_2_28;
wire n_0_329;
wire n_0_2_29;
wire n_0_394;
wire n_0_2_30;
wire n_0_330;
wire n_0_2_31;
wire n_0_395;
wire n_0_2_32;
wire n_0_331;
wire n_0_2_33;
wire n_0_396;
wire n_0_2_34;
wire n_0_332;
wire n_0_2_35;
wire n_0_397;
wire n_0_2_36;
wire n_0_333;
wire n_0_2_37;
wire n_0_398;
wire n_0_2_38;
wire n_0_334;
wire n_0_2_39;
wire n_0_399;
wire n_0_2_40;
wire n_0_335;
wire n_0_2_41;
wire n_0_400;
wire n_0_2_42;
wire n_0_336;
wire n_0_2_43;
wire n_0_401;
wire n_0_2_44;
wire n_0_337;
wire n_0_2_45;
wire n_0_402;
wire n_0_2_46;
wire n_0_338;
wire n_0_2_47;
wire n_0_403;
wire n_0_2_48;
wire n_0_339;
wire n_0_2_49;
wire n_0_404;
wire n_0_2_50;
wire n_0_340;
wire n_0_2_51;
wire n_0_405;
wire n_0_2_52;
wire n_0_341;
wire n_0_2_53;
wire n_0_406;
wire n_0_2_54;
wire n_0_342;
wire n_0_2_55;
wire n_0_407;
wire n_0_2_56;
wire n_0_343;
wire n_0_2_57;
wire n_0_408;
wire n_0_2_58;
wire n_0_344;
wire n_0_2_59;
wire n_0_409;
wire n_0_2_60;
wire n_0_345;
wire n_0_2_61;
wire n_0_410;
wire n_0_2_62;
wire n_0_346;
wire n_0_2_63;
wire n_0_411;
wire n_0_2_64;
wire n_0_347;
wire n_0_2_65;
wire n_0_412;
wire n_0_2_66;
wire n_0_348;
wire n_0_2_67;
wire n_0_413;
wire n_0_2_68;
wire n_0_349;
wire n_0_2_69;
wire n_0_414;
wire n_0_2_70;
wire n_0_350;
wire n_0_2_71;
wire n_0_415;
wire n_0_2_72;
wire n_0_351;
wire n_0_2_73;
wire n_0_416;
wire n_0_2_74;
wire n_0_352;
wire n_0_2_75;
wire n_0_417;
wire n_0_2_76;
wire n_0_353;
wire n_0_2_77;
wire n_0_418;
wire n_0_2_78;
wire n_0_354;
wire n_0_2_79;
wire n_0_419;
wire n_0_2_80;
wire n_0_355;
wire n_0_2_81;
wire n_0_420;
wire n_0_2_82;
wire n_0_356;
wire n_0_2_83;
wire n_0_421;
wire n_0_2_84;
wire n_0_357;
wire n_0_2_85;
wire n_0_422;
wire n_0_2_86;
wire n_0_358;
wire n_0_2_87;
wire n_0_423;
wire n_0_2_88;
wire n_0_359;
wire n_0_2_89;
wire n_0_424;
wire n_0_2_90;
wire n_0_360;
wire n_0_2_91;
wire n_0_425;
wire n_0_2_92;
wire n_0_361;
wire n_0_2_93;
wire n_0_426;
wire n_0_2_94;
wire n_0_362;
wire n_0_2_95;
wire n_0_427;
wire n_0_2_96;
wire n_0_363;
wire n_0_2_97;
wire n_0_428;
wire n_0_2_98;
wire n_0_364;
wire n_0_2_99;
wire n_0_429;
wire n_0_2_100;
wire n_0_365;
wire n_0_2_101;
wire n_0_430;
wire n_0_2_102;
wire n_0_366;
wire n_0_2_103;
wire n_0_431;
wire n_0_2_104;
wire n_0_367;
wire n_0_2_105;
wire n_0_432;
wire n_0_2_106;
wire n_0_368;
wire n_0_2_107;
wire n_0_433;
wire n_0_2_108;
wire n_0_369;
wire n_0_2_109;
wire n_0_434;
wire n_0_2_110;
wire n_0_370;
wire n_0_2_111;
wire n_0_435;
wire n_0_2_112;
wire n_0_371;
wire n_0_2_113;
wire n_0_436;
wire n_0_2_114;
wire n_0_372;
wire n_0_2_115;
wire n_0_437;
wire n_0_2_116;
wire n_0_373;
wire n_0_2_117;
wire n_0_438;
wire n_0_2_118;
wire n_0_374;
wire n_0_2_119;
wire n_0_439;
wire n_0_2_120;
wire n_0_375;
wire n_0_2_121;
wire n_0_440;
wire n_0_2_122;
wire n_0_376;
wire n_0_2_123;
wire n_0_441;
wire n_0_2_124;
wire n_0_377;
wire n_0_2_125;
wire n_0_442;
wire n_0_2_126;
wire n_0_378;
wire n_0_2_127;
wire n_0_443;
wire n_0_2_128;
wire n_0_379;
wire n_0_2_129;
wire n_0_444;
wire n_0_2_130;
wire n_0_380;
wire n_0_2_131;
wire n_0_445;
wire n_0_2_132;
wire n_0_381;
wire n_0_2_133;
wire n_0_446;
wire n_0_2_134;
wire n_0_382;
wire n_0_2_135;
wire n_0_447;
wire n_0_2_136;
wire n_0_383;
wire n_0_2_137;
wire n_0_448;
wire n_0_2_138;
wire n_0_384;
wire n_0_2_139;
wire n_0_449;
wire n_0_2_140;
wire n_0_385;
wire n_0_2_141;
wire n_0_450;
wire n_0_2_142;
wire n_0_386;
wire n_0_2_143;
wire n_0_451;
wire n_0_2_144;
wire n_0_387;
wire n_0_2_145;
wire n_0_452;
wire n_0_2_146;
wire n_0_388;
wire n_0_2_147;
wire n_0_2_148;
wire n_0_2_149;
wire n_0_2_150;
wire n_0_2_151;
wire n_0_2_152;
wire n_0_2_153;
wire n_0_2_154;
wire n_0_2_155;
wire n_0_2_156;
wire n_0_2_157;
wire n_0_2_158;
wire n_0_2_159;
wire n_0_2_160;
wire n_0_2_161;
wire n_0_2_162;
wire n_0_2_163;
wire n_0_2_164;
wire n_0_2_165;
wire n_0_2_166;
wire n_0_2_167;
wire n_0_2_168;
wire n_0_2_169;
wire n_0_2_170;
wire n_0_2_171;
wire n_0_2_172;
wire n_0_2_173;
wire n_0_2_174;
wire n_0_2_175;
wire n_0_2_176;
wire n_0_2_177;
wire n_0_2_178;
wire n_0_2_179;
wire n_0_389;
wire n_0_2_180;
wire n_0_2_181;
wire n_0_2_182;
wire n_0_2_183;
wire n_0_260;
wire n_0_2_184;
wire n_0_2_185;
wire n_0_261;
wire n_0_2_186;
wire n_0_2_187;
wire n_0_2_188;
wire n_0_262;
wire n_0_2_189;
wire n_0_263;
wire n_0_2_190;
wire n_0_2_191;
wire n_0_2_192;
wire n_0_2_193;
wire n_0_2_194;
wire n_0_264;
wire n_0_2_195;
wire n_0_2_196;
wire n_0_2_197;
wire n_0_265;
wire n_0_2_198;
wire n_0_2_199;
wire n_0_2_200;
wire n_0_2_201;
wire n_0_2_202;
wire n_0_266;
wire n_0_2_203;
wire n_0_2_204;
wire n_0_2_205;
wire n_0_2_206;
wire n_0_267;
wire n_0_2_207;
wire n_0_2_208;
wire n_0_2_209;
wire n_0_2_210;
wire n_0_2_211;
wire n_0_268;
wire n_0_2_212;
wire n_0_2_213;
wire n_0_2_214;
wire n_0_2_215;
wire n_0_269;
wire n_0_2_216;
wire n_0_2_217;
wire n_0_2_218;
wire n_0_2_219;
wire n_0_2_220;
wire n_0_2_221;
wire n_0_2_222;
wire n_0_2_223;
wire n_0_270;
wire n_0_2_224;
wire n_0_2_225;
wire n_0_2_226;
wire n_0_2_227;
wire n_0_2_228;
wire n_0_2_229;
wire n_0_271;
wire n_0_2_230;
wire n_0_2_231;
wire n_0_2_232;
wire n_0_272;
wire n_0_2_233;
wire n_0_2_234;
wire n_0_2_235;
wire n_0_273;
wire n_0_2_236;
wire n_0_2_237;
wire n_0_2_238;
wire n_0_274;
wire n_0_2_239;
wire n_0_2_240;
wire n_0_2_241;
wire n_0_275;
wire n_0_2_242;
wire n_0_2_243;
wire n_0_2_244;
wire n_0_2_245;
wire n_0_2_246;
wire n_0_2_247;
wire n_0_2_248;
wire n_0_276;
wire n_0_2_249;
wire n_0_2_250;
wire n_0_2_251;
wire n_0_2_252;
wire n_0_2_253;
wire n_0_2_254;
wire n_0_277;
wire n_0_2_255;
wire n_0_2_256;
wire n_0_2_257;
wire n_0_2_258;
wire n_0_2_259;
wire n_0_278;
wire n_0_2_260;
wire n_0_2_261;
wire n_0_2_262;
wire n_0_2_263;
wire n_0_2_264;
wire n_0_279;
wire n_0_2_265;
wire n_0_2_266;
wire n_0_2_267;
wire n_0_2_268;
wire n_0_2_269;
wire n_0_2_270;
wire n_0_2_271;
wire n_0_280;
wire n_0_2_272;
wire n_0_2_273;
wire n_0_2_274;
wire n_0_2_275;
wire n_0_2_276;
wire n_0_2_277;
wire n_0_281;
wire n_0_2_278;
wire n_0_2_279;
wire n_0_2_280;
wire n_0_2_281;
wire n_0_2_282;
wire n_0_2_283;
wire n_0_282;
wire n_0_2_284;
wire n_0_2_285;
wire n_0_2_286;
wire n_0_2_287;
wire n_0_2_288;
wire n_0_2_289;
wire n_0_283;
wire n_0_2_290;
wire n_0_2_291;
wire n_0_2_292;
wire n_0_2_293;
wire n_0_2_294;
wire n_0_2_295;
wire n_0_2_296;
wire n_0_2_297;
wire n_0_284;
wire n_0_2_298;
wire n_0_2_299;
wire n_0_2_300;
wire n_0_2_301;
wire n_0_2_302;
wire n_0_2_303;
wire n_0_2_304;
wire n_0_285;
wire n_0_2_305;
wire n_0_2_306;
wire n_0_2_307;
wire n_0_2_308;
wire n_0_2_309;
wire n_0_2_310;
wire n_0_286;
wire n_0_2_311;
wire n_0_2_312;
wire n_0_2_313;
wire n_0_2_314;
wire n_0_2_315;
wire n_0_2_316;
wire n_0_2_317;
wire n_0_287;
wire n_0_2_318;
wire n_0_2_319;
wire n_0_2_320;
wire n_0_2_321;
wire n_0_2_322;
wire n_0_2_323;
wire n_0_2_324;
wire n_0_288;
wire n_0_2_325;
wire n_0_2_326;
wire n_0_2_327;
wire n_0_2_328;
wire n_0_2_329;
wire n_0_2_330;
wire n_0_2_331;
wire n_0_289;
wire n_0_2_332;
wire n_0_2_333;
wire n_0_2_334;
wire n_0_2_335;
wire n_0_2_336;
wire n_0_2_337;
wire n_0_2_338;
wire n_0_290;
wire n_0_2_339;
wire n_0_2_340;
wire n_0_2_341;
wire n_0_2_342;
wire n_0_2_343;
wire n_0_2_344;
wire n_0_2_345;
wire n_0_291;
wire n_0_2_346;
wire n_0_2_347;
wire n_0_2_348;
wire n_0_2_349;
wire n_0_2_350;
wire n_0_292;
wire n_0_2_351;
wire n_0_2_352;
wire n_0_2_353;
wire n_0_2_354;
wire n_0_293;
wire n_0_2_355;
wire n_0_2_356;
wire n_0_2_357;
wire n_0_2_358;
wire n_0_294;
wire n_0_2_359;
wire n_0_2_360;
wire n_0_2_361;
wire n_0_2_362;
wire n_0_295;
wire n_0_2_363;
wire n_0_2_364;
wire n_0_2_365;
wire n_0_2_366;
wire n_0_296;
wire n_0_2_367;
wire n_0_2_368;
wire n_0_2_369;
wire n_0_2_370;
wire n_0_297;
wire n_0_2_371;
wire n_0_2_372;
wire n_0_2_373;
wire n_0_2_374;
wire n_0_298;
wire n_0_2_375;
wire n_0_2_376;
wire n_0_2_377;
wire n_0_2_378;
wire n_0_299;
wire n_0_2_379;
wire n_0_2_380;
wire n_0_2_381;
wire n_0_2_382;
wire n_0_2_383;
wire n_0_300;
wire n_0_2_384;
wire n_0_2_385;
wire n_0_2_386;
wire n_0_2_387;
wire n_0_2_388;
wire n_0_301;
wire n_0_2_389;
wire n_0_2_390;
wire n_0_2_391;
wire n_0_2_392;
wire n_0_302;
wire n_0_2_393;
wire n_0_2_394;
wire n_0_2_395;
wire n_0_2_396;
wire n_0_2_397;
wire n_0_303;
wire n_0_2_398;
wire n_0_2_399;
wire n_0_2_400;
wire n_0_2_401;
wire n_0_2_402;
wire n_0_304;
wire n_0_2_403;
wire n_0_2_404;
wire n_0_2_405;
wire n_0_2_406;
wire n_0_2_407;
wire n_0_305;
wire n_0_2_408;
wire n_0_2_409;
wire n_0_2_410;
wire n_0_2_411;
wire n_0_2_412;
wire n_0_306;
wire n_0_2_413;
wire n_0_2_414;
wire n_0_2_415;
wire n_0_2_416;
wire n_0_2_417;
wire n_0_307;
wire n_0_2_418;
wire n_0_2_419;
wire n_0_2_420;
wire n_0_2_421;
wire n_0_2_422;
wire n_0_308;
wire n_0_2_423;
wire n_0_2_424;
wire n_0_2_425;
wire n_0_309;
wire n_0_2_426;
wire n_0_2_427;
wire n_0_2_428;
wire n_0_310;
wire n_0_2_429;
wire n_0_2_430;
wire n_0_2_431;
wire n_0_311;
wire n_0_2_432;
wire n_0_2_433;
wire n_0_2_434;
wire n_0_312;
wire n_0_2_435;
wire n_0_2_436;
wire n_0_2_437;
wire n_0_313;
wire n_0_2_438;
wire n_0_2_439;
wire n_0_2_440;
wire n_0_314;
wire n_0_2_441;
wire n_0_2_442;
wire n_0_2_443;
wire n_0_315;
wire n_0_2_444;
wire n_0_2_445;
wire n_0_2_446;
wire n_0_2_447;
wire n_0_2_448;
wire n_0_316;
wire n_0_2_449;
wire n_0_2_450;
wire n_0_2_451;
wire n_0_2_452;
wire n_0_317;
wire n_0_2_453;
wire n_0_2_454;
wire n_0_2_455;
wire n_0_2_456;
wire n_0_318;
wire n_0_2_457;
wire n_0_2_458;
wire n_0_2_459;
wire n_0_2_460;
wire n_0_319;
wire n_0_2_461;
wire n_0_2_462;
wire n_0_320;
wire n_0_2_463;
wire n_0_2_464;
wire n_0_321;
wire n_0_2_465;
wire n_0_2_466;
wire n_0_2_467;
wire n_0_2_468;
wire n_0_2_469;
wire n_0_322;
wire n_0_2_470;
wire n_0_2_471;
wire n_0_2_472;
wire n_0_323;
wire \outmultiplicand_reg[31] ;
wire \outmultiplicand_reg[30] ;
wire \outmultiplicand_reg[29] ;
wire \outmultiplicand_reg[28] ;
wire \outmultiplicand_reg[27] ;
wire \outmultiplicand_reg[26] ;
wire \outmultiplicand_reg[25] ;
wire \outmultiplicand_reg[24] ;
wire \outmultiplicand_reg[23] ;
wire \outmultiplicand_reg[22] ;
wire \outmultiplicand_reg[21] ;
wire \outmultiplicand_reg[20] ;
wire \outmultiplicand_reg[19] ;
wire \outmultiplicand_reg[18] ;
wire \outmultiplicand_reg[17] ;
wire \outmultiplicand_reg[16] ;
wire \outmultiplicand_reg[15] ;
wire \outmultiplicand_reg[14] ;
wire \outmultiplicand_reg[13] ;
wire \outmultiplicand_reg[12] ;
wire \outmultiplicand_reg[11] ;
wire \outmultiplicand_reg[10] ;
wire \outmultiplicand_reg[9] ;
wire \outmultiplicand_reg[8] ;
wire \outmultiplicand_reg[7] ;
wire \outmultiplicand_reg[6] ;
wire \outmultiplicand_reg[5] ;
wire \outmultiplicand_reg[4] ;
wire \outmultiplicand_reg[3] ;
wire \outmultiplicand_reg[2] ;
wire \outmultiplicand_reg[1] ;
wire \outmultiplicand_reg[0] ;
wire n_0_0;
wire \accumulator[63] ;
wire \accumulator[62] ;
wire \accumulator[61] ;
wire \accumulator[60] ;
wire \accumulator[59] ;
wire \accumulator[58] ;
wire \accumulator[57] ;
wire \accumulator[56] ;
wire \accumulator[55] ;
wire \accumulator[54] ;
wire \accumulator[53] ;
wire \accumulator[52] ;
wire \accumulator[51] ;
wire \accumulator[50] ;
wire \accumulator[49] ;
wire \accumulator[48] ;
wire \accumulator[47] ;
wire \accumulator[46] ;
wire \accumulator[45] ;
wire \accumulator[44] ;
wire \accumulator[43] ;
wire \accumulator[42] ;
wire \accumulator[41] ;
wire \accumulator[40] ;
wire \accumulator[39] ;
wire \accumulator[38] ;
wire \accumulator[37] ;
wire \accumulator[36] ;
wire \accumulator[35] ;
wire \accumulator[34] ;
wire \accumulator[33] ;
wire \accumulator[32] ;
wire \accumulator[31] ;
wire \accumulator[30] ;
wire \accumulator[29] ;
wire \accumulator[28] ;
wire \accumulator[27] ;
wire \accumulator[26] ;
wire \accumulator[25] ;
wire \accumulator[24] ;
wire \accumulator[23] ;
wire \accumulator[22] ;
wire \accumulator[21] ;
wire \accumulator[20] ;
wire \accumulator[19] ;
wire \accumulator[18] ;
wire \accumulator[17] ;
wire \accumulator[16] ;
wire \accumulator[15] ;
wire \accumulator[14] ;
wire \accumulator[13] ;
wire \accumulator[12] ;
wire \accumulator[11] ;
wire \accumulator[10] ;
wire \accumulator[9] ;
wire \accumulator[8] ;
wire \accumulator[7] ;
wire \accumulator[6] ;
wire \accumulator[5] ;
wire \accumulator[4] ;
wire \accumulator[3] ;
wire \accumulator[2] ;
wire \accumulator[1] ;
wire \accumulator[0] ;
wire \multiplier1[31] ;
wire \multiplier1[30] ;
wire \multiplier1[29] ;
wire \multiplier1[28] ;
wire \multiplier1[27] ;
wire \multiplier1[26] ;
wire \multiplier1[25] ;
wire \multiplier1[24] ;
wire \multiplier1[23] ;
wire \multiplier1[22] ;
wire \multiplier1[21] ;
wire \multiplier1[20] ;
wire \multiplier1[19] ;
wire \multiplier1[18] ;
wire \multiplier1[17] ;
wire \multiplier1[16] ;
wire \multiplier1[15] ;
wire \multiplier1[14] ;
wire \multiplier1[13] ;
wire \multiplier1[12] ;
wire \multiplier1[11] ;
wire \multiplier1[10] ;
wire \multiplier1[9] ;
wire \multiplier1[8] ;
wire \multiplier1[7] ;
wire \multiplier1[6] ;
wire \multiplier1[5] ;
wire \multiplier1[4] ;
wire \multiplier1[3] ;
wire \multiplier1[2] ;
wire \multiplier1[1] ;
wire \multiplier1[0] ;
wire \counter[5] ;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire spw__n338;
wire spw__n337;
wire spw__n326;
wire spw__n325;
wire spw__n324;
wire spw__n323;
wire spw__n312;
wire spw__n311;
wire spw__n310;
wire spw__n309;
wire spw__n156;
wire spw__n155;
wire spw__n125;
wire spw__n124;
wire spw__n123;
wire spt__n28;
wire spt__n25;
wire spc__n22;
wire spc__n19;
wire spc__n16;
wire sps__n13;
wire sps__n10;
wire sps__n7;
wire sps__n4;
wire sps__n1;
wire \multiplicand1[31] ;
wire \multiplicand1[30] ;
wire \multiplicand1[29] ;
wire \multiplicand1[28] ;
wire \multiplicand1[27] ;
wire \multiplicand1[26] ;
wire \multiplicand1[25] ;
wire \multiplicand1[24] ;
wire \multiplicand1[23] ;
wire \multiplicand1[22] ;
wire \multiplicand1[21] ;
wire \multiplicand1[20] ;
wire \multiplicand1[19] ;
wire \multiplicand1[18] ;
wire \multiplicand1[17] ;
wire \multiplicand1[16] ;
wire \multiplicand1[15] ;
wire \multiplicand1[14] ;
wire \multiplicand1[13] ;
wire \multiplicand1[12] ;
wire \multiplicand1[11] ;
wire \multiplicand1[10] ;
wire \multiplicand1[9] ;
wire \multiplicand1[8] ;
wire \multiplicand1[7] ;
wire \multiplicand1[6] ;
wire \multiplicand1[5] ;
wire \multiplicand1[4] ;
wire \multiplicand1[3] ;
wire \multiplicand1[2] ;
wire \multiplicand1[1] ;
wire \multiplicand1[0] ;
wire negative_product_flag;
wire n_0_1;
wire n_0_228;
wire uc_0;
wire uc_1;
wire uc_2;


CLKGATETST_X1 clk_gate_negative_product_flag_reg (.GCK (n_0_228), .CK (clk), .E (set_signal), .SE (1'b0 ));
CLKGATETST_X1 clk_gate_outmultiplicand_reg_reg (.GCK (n_0_1), .CK (clk), .E (n_0_453), .SE (1'b0 ));
DFF_X1 negative_product_flag_reg (.Q (negative_product_flag), .CK (n_0_228), .D (n_0_191));
DFF_X1 \multiplicand1_reg[0]  (.Q (\multiplicand1[0] ), .CK (n_0_228), .D (\multiplicand_reg[0] ));
DFF_X1 \multiplicand1_reg[1]  (.Q (\multiplicand1[1] ), .CK (n_0_228), .D (n_0_192));
DFF_X1 \multiplicand1_reg[2]  (.Q (\multiplicand1[2] ), .CK (n_0_228), .D (n_0_193));
DFF_X1 \multiplicand1_reg[3]  (.Q (\multiplicand1[3] ), .CK (n_0_228), .D (n_0_194));
DFF_X1 \multiplicand1_reg[4]  (.Q (\multiplicand1[4] ), .CK (n_0_228), .D (n_0_195));
DFF_X1 \multiplicand1_reg[5]  (.Q (\multiplicand1[5] ), .CK (n_0_228), .D (n_0_196));
DFF_X1 \multiplicand1_reg[6]  (.Q (\multiplicand1[6] ), .CK (n_0_228), .D (n_0_197));
DFF_X1 \multiplicand1_reg[7]  (.Q (\multiplicand1[7] ), .CK (n_0_228), .D (n_0_198));
DFF_X1 \multiplicand1_reg[8]  (.Q (\multiplicand1[8] ), .CK (n_0_228), .D (n_0_199));
DFF_X1 \multiplicand1_reg[9]  (.Q (\multiplicand1[9] ), .CK (n_0_228), .D (n_0_200));
DFF_X1 \multiplicand1_reg[10]  (.Q (\multiplicand1[10] ), .CK (n_0_228), .D (n_0_201));
DFF_X1 \multiplicand1_reg[11]  (.Q (\multiplicand1[11] ), .CK (n_0_228), .D (n_0_202));
DFF_X1 \multiplicand1_reg[12]  (.Q (\multiplicand1[12] ), .CK (n_0_228), .D (n_0_203));
DFF_X1 \multiplicand1_reg[13]  (.Q (\multiplicand1[13] ), .CK (n_0_228), .D (n_0_204));
DFF_X1 \multiplicand1_reg[14]  (.Q (\multiplicand1[14] ), .CK (n_0_228), .D (n_0_205));
DFF_X1 \multiplicand1_reg[15]  (.Q (\multiplicand1[15] ), .CK (n_0_228), .D (n_0_206));
DFF_X1 \multiplicand1_reg[16]  (.Q (\multiplicand1[16] ), .CK (n_0_228), .D (n_0_207));
DFF_X1 \multiplicand1_reg[17]  (.Q (\multiplicand1[17] ), .CK (n_0_228), .D (n_0_208));
DFF_X1 \multiplicand1_reg[18]  (.Q (\multiplicand1[18] ), .CK (n_0_228), .D (n_0_209));
DFF_X1 \multiplicand1_reg[19]  (.Q (\multiplicand1[19] ), .CK (n_0_228), .D (n_0_210));
DFF_X1 \multiplicand1_reg[20]  (.Q (\multiplicand1[20] ), .CK (n_0_228), .D (n_0_211));
DFF_X1 \multiplicand1_reg[21]  (.Q (\multiplicand1[21] ), .CK (n_0_228), .D (n_0_212));
DFF_X1 \multiplicand1_reg[22]  (.Q (\multiplicand1[22] ), .CK (n_0_228), .D (n_0_213));
DFF_X1 \multiplicand1_reg[23]  (.Q (\multiplicand1[23] ), .CK (n_0_228), .D (n_0_214));
DFF_X1 \multiplicand1_reg[24]  (.Q (\multiplicand1[24] ), .CK (n_0_228), .D (n_0_215));
DFF_X1 \multiplicand1_reg[25]  (.Q (\multiplicand1[25] ), .CK (n_0_228), .D (n_0_216));
DFF_X1 \multiplicand1_reg[26]  (.Q (\multiplicand1[26] ), .CK (n_0_228), .D (n_0_217));
DFF_X1 \multiplicand1_reg[27]  (.Q (\multiplicand1[27] ), .CK (n_0_228), .D (n_0_218));
DFF_X1 \multiplicand1_reg[28]  (.Q (\multiplicand1[28] ), .CK (n_0_228), .D (n_0_219));
DFF_X1 \multiplicand1_reg[29]  (.Q (\multiplicand1[29] ), .CK (n_0_228), .D (n_0_220));
DFF_X1 \multiplicand1_reg[30]  (.Q (\multiplicand1[30] ), .CK (n_0_228), .D (n_0_221));
DFF_X1 \multiplicand1_reg[31]  (.Q (\multiplicand1[31] ), .CK (n_0_228), .D (n_0_222));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (clk), .D (n_0_255));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (clk), .D (n_0_256));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (clk), .D (n_0_257));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (clk), .D (n_0_258));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (clk), .D (n_0_259));
DFF_X1 \counter_reg[5]  (.Q (\counter[5] ), .CK (clk), .D (n_0_324));
DFF_X1 \multiplier1_reg[0]  (.Q (\multiplier1[0] ), .CK (n_0_228), .D (\multiplier_reg[0] ));
DFF_X1 \multiplier1_reg[1]  (.Q (\multiplier1[1] ), .CK (n_0_228), .D (n_0_223));
DFF_X1 \multiplier1_reg[2]  (.Q (\multiplier1[2] ), .CK (n_0_228), .D (n_0_224));
DFF_X1 \multiplier1_reg[3]  (.Q (\multiplier1[3] ), .CK (n_0_228), .D (n_0_225));
DFF_X1 \multiplier1_reg[4]  (.Q (\multiplier1[4] ), .CK (n_0_228), .D (n_0_226));
DFF_X1 \multiplier1_reg[5]  (.Q (\multiplier1[5] ), .CK (n_0_228), .D (n_0_227));
DFF_X1 \multiplier1_reg[6]  (.Q (\multiplier1[6] ), .CK (n_0_228), .D (n_0_229));
DFF_X1 \multiplier1_reg[7]  (.Q (\multiplier1[7] ), .CK (n_0_228), .D (n_0_230));
DFF_X1 \multiplier1_reg[8]  (.Q (\multiplier1[8] ), .CK (n_0_228), .D (n_0_231));
DFF_X1 \multiplier1_reg[9]  (.Q (\multiplier1[9] ), .CK (n_0_228), .D (n_0_232));
DFF_X1 \multiplier1_reg[10]  (.Q (\multiplier1[10] ), .CK (n_0_228), .D (n_0_233));
DFF_X1 \multiplier1_reg[11]  (.Q (\multiplier1[11] ), .CK (n_0_228), .D (n_0_234));
DFF_X1 \multiplier1_reg[12]  (.Q (\multiplier1[12] ), .CK (n_0_228), .D (n_0_235));
DFF_X1 \multiplier1_reg[13]  (.Q (\multiplier1[13] ), .CK (n_0_228), .D (n_0_236));
DFF_X1 \multiplier1_reg[14]  (.Q (\multiplier1[14] ), .CK (n_0_228), .D (n_0_237));
DFF_X1 \multiplier1_reg[15]  (.Q (\multiplier1[15] ), .CK (n_0_228), .D (n_0_238));
DFF_X1 \multiplier1_reg[16]  (.Q (\multiplier1[16] ), .CK (n_0_228), .D (n_0_239));
DFF_X1 \multiplier1_reg[17]  (.Q (\multiplier1[17] ), .CK (n_0_228), .D (n_0_240));
DFF_X1 \multiplier1_reg[18]  (.Q (\multiplier1[18] ), .CK (n_0_228), .D (n_0_241));
DFF_X1 \multiplier1_reg[19]  (.Q (\multiplier1[19] ), .CK (n_0_228), .D (n_0_242));
DFF_X1 \multiplier1_reg[20]  (.Q (\multiplier1[20] ), .CK (n_0_228), .D (n_0_243));
DFF_X1 \multiplier1_reg[21]  (.Q (\multiplier1[21] ), .CK (n_0_228), .D (n_0_244));
DFF_X1 \multiplier1_reg[22]  (.Q (\multiplier1[22] ), .CK (n_0_228), .D (n_0_245));
DFF_X1 \multiplier1_reg[23]  (.Q (\multiplier1[23] ), .CK (n_0_228), .D (n_0_246));
DFF_X1 \multiplier1_reg[24]  (.Q (\multiplier1[24] ), .CK (n_0_228), .D (n_0_247));
DFF_X1 \multiplier1_reg[25]  (.Q (\multiplier1[25] ), .CK (n_0_228), .D (n_0_248));
DFF_X1 \multiplier1_reg[26]  (.Q (\multiplier1[26] ), .CK (n_0_228), .D (n_0_249));
DFF_X1 \multiplier1_reg[27]  (.Q (\multiplier1[27] ), .CK (n_0_228), .D (n_0_250));
DFF_X1 \multiplier1_reg[28]  (.Q (\multiplier1[28] ), .CK (n_0_228), .D (n_0_251));
DFF_X1 \multiplier1_reg[29]  (.Q (\multiplier1[29] ), .CK (n_0_228), .D (n_0_252));
DFF_X1 \multiplier1_reg[30]  (.Q (\multiplier1[30] ), .CK (n_0_228), .D (n_0_253));
DFF_X1 \multiplier1_reg[31]  (.Q (\multiplier1[31] ), .CK (n_0_228), .D (n_0_254));
DFF_X1 \accumulator_reg[0]  (.Q (spw__n125), .CK (n_0_0), .D (n_0_325));
DFF_X1 \accumulator_reg[1]  (.Q (\accumulator[1] ), .CK (n_0_0), .D (n_0_326));
DFF_X1 \accumulator_reg[2]  (.Q (\accumulator[2] ), .CK (n_0_0), .D (n_0_327));
DFF_X1 \accumulator_reg[3]  (.Q (\accumulator[3] ), .CK (n_0_0), .D (n_0_328));
DFF_X1 \accumulator_reg[4]  (.Q (\accumulator[4] ), .CK (n_0_0), .D (n_0_329));
DFF_X1 \accumulator_reg[5]  (.Q (\accumulator[5] ), .CK (n_0_0), .D (n_0_330));
DFF_X1 \accumulator_reg[6]  (.Q (\accumulator[6] ), .CK (n_0_0), .D (n_0_331));
DFF_X1 \accumulator_reg[7]  (.Q (\accumulator[7] ), .CK (n_0_0), .D (n_0_332));
DFF_X1 \accumulator_reg[8]  (.Q (\accumulator[8] ), .CK (n_0_0), .D (n_0_333));
DFF_X1 \accumulator_reg[9]  (.Q (\accumulator[9] ), .CK (n_0_0), .D (n_0_334));
DFF_X1 \accumulator_reg[10]  (.Q (\accumulator[10] ), .CK (n_0_0), .D (n_0_335));
DFF_X1 \accumulator_reg[11]  (.Q (\accumulator[11] ), .CK (n_0_0), .D (n_0_336));
DFF_X1 \accumulator_reg[12]  (.Q (\accumulator[12] ), .CK (n_0_0), .D (n_0_337));
DFF_X1 \accumulator_reg[13]  (.Q (\accumulator[13] ), .CK (n_0_0), .D (n_0_338));
DFF_X1 \accumulator_reg[14]  (.Q (\accumulator[14] ), .CK (n_0_0), .D (n_0_339));
DFF_X1 \accumulator_reg[15]  (.Q (\accumulator[15] ), .CK (n_0_0), .D (n_0_340));
DFF_X1 \accumulator_reg[16]  (.Q (\accumulator[16] ), .CK (n_0_0), .D (n_0_341));
DFF_X1 \accumulator_reg[17]  (.Q (\accumulator[17] ), .CK (n_0_0), .D (n_0_342));
DFF_X1 \accumulator_reg[18]  (.Q (\accumulator[18] ), .CK (n_0_0), .D (n_0_343));
DFF_X1 \accumulator_reg[19]  (.Q (\accumulator[19] ), .CK (n_0_0), .D (n_0_344));
DFF_X1 \accumulator_reg[20]  (.Q (\accumulator[20] ), .CK (n_0_0), .D (n_0_345));
DFF_X1 \accumulator_reg[21]  (.Q (\accumulator[21] ), .CK (n_0_0), .D (n_0_346));
DFF_X1 \accumulator_reg[22]  (.Q (\accumulator[22] ), .CK (n_0_0), .D (n_0_347));
DFF_X1 \accumulator_reg[23]  (.Q (\accumulator[23] ), .CK (n_0_0), .D (n_0_348));
DFF_X1 \accumulator_reg[24]  (.Q (\accumulator[24] ), .CK (n_0_0), .D (n_0_349));
DFF_X1 \accumulator_reg[25]  (.Q (\accumulator[25] ), .CK (n_0_0), .D (n_0_350));
DFF_X1 \accumulator_reg[26]  (.Q (\accumulator[26] ), .CK (n_0_0), .D (n_0_351));
DFF_X1 \accumulator_reg[27]  (.Q (\accumulator[27] ), .CK (n_0_0), .D (n_0_352));
DFF_X1 \accumulator_reg[28]  (.Q (\accumulator[28] ), .CK (n_0_0), .D (n_0_353));
DFF_X1 \accumulator_reg[29]  (.Q (\accumulator[29] ), .CK (n_0_0), .D (n_0_354));
DFF_X1 \accumulator_reg[30]  (.Q (\accumulator[30] ), .CK (n_0_0), .D (n_0_355));
DFF_X1 \accumulator_reg[31]  (.Q (\accumulator[31] ), .CK (n_0_0), .D (n_0_356));
DFF_X1 \accumulator_reg[32]  (.Q (\accumulator[32] ), .CK (n_0_0), .D (n_0_357));
DFF_X1 \accumulator_reg[33]  (.Q (\accumulator[33] ), .CK (n_0_0), .D (n_0_358));
DFF_X1 \accumulator_reg[34]  (.Q (\accumulator[34] ), .CK (n_0_0), .D (n_0_359));
DFF_X1 \accumulator_reg[35]  (.Q (\accumulator[35] ), .CK (n_0_0), .D (n_0_360));
DFF_X1 \accumulator_reg[36]  (.Q (\accumulator[36] ), .CK (n_0_0), .D (n_0_361));
DFF_X1 \accumulator_reg[37]  (.Q (\accumulator[37] ), .CK (n_0_0), .D (n_0_362));
DFF_X1 \accumulator_reg[38]  (.Q (\accumulator[38] ), .CK (n_0_0), .D (n_0_363));
DFF_X1 \accumulator_reg[39]  (.Q (\accumulator[39] ), .CK (n_0_0), .D (n_0_364));
DFF_X1 \accumulator_reg[40]  (.Q (\accumulator[40] ), .CK (n_0_0), .D (n_0_365));
DFF_X1 \accumulator_reg[41]  (.Q (\accumulator[41] ), .CK (n_0_0), .D (n_0_366));
DFF_X1 \accumulator_reg[42]  (.Q (\accumulator[42] ), .CK (n_0_0), .D (n_0_367));
DFF_X1 \accumulator_reg[43]  (.Q (\accumulator[43] ), .CK (n_0_0), .D (n_0_368));
DFF_X1 \accumulator_reg[44]  (.Q (\accumulator[44] ), .CK (n_0_0), .D (n_0_369));
DFF_X1 \accumulator_reg[45]  (.Q (\accumulator[45] ), .CK (n_0_0), .D (n_0_370));
DFF_X1 \accumulator_reg[46]  (.Q (\accumulator[46] ), .CK (n_0_0), .D (n_0_371));
DFF_X1 \accumulator_reg[47]  (.Q (\accumulator[47] ), .CK (n_0_0), .D (n_0_372));
DFF_X1 \accumulator_reg[48]  (.Q (\accumulator[48] ), .CK (n_0_0), .D (n_0_373));
DFF_X1 \accumulator_reg[49]  (.Q (\accumulator[49] ), .CK (n_0_0), .D (n_0_374));
DFF_X1 \accumulator_reg[50]  (.Q (\accumulator[50] ), .CK (n_0_0), .D (n_0_375));
DFF_X1 \accumulator_reg[51]  (.Q (\accumulator[51] ), .CK (n_0_0), .D (n_0_376));
DFF_X1 \accumulator_reg[52]  (.Q (\accumulator[52] ), .CK (n_0_0), .D (n_0_377));
DFF_X1 \accumulator_reg[53]  (.Q (\accumulator[53] ), .CK (n_0_0), .D (n_0_378));
DFF_X1 \accumulator_reg[54]  (.Q (\accumulator[54] ), .CK (n_0_0), .D (n_0_379));
DFF_X1 \accumulator_reg[55]  (.Q (\accumulator[55] ), .CK (n_0_0), .D (n_0_380));
DFF_X1 \accumulator_reg[56]  (.Q (\accumulator[56] ), .CK (n_0_0), .D (n_0_381));
DFF_X1 \accumulator_reg[57]  (.Q (\accumulator[57] ), .CK (n_0_0), .D (n_0_382));
DFF_X1 \accumulator_reg[58]  (.Q (\accumulator[58] ), .CK (n_0_0), .D (n_0_383));
DFF_X1 \accumulator_reg[59]  (.Q (\accumulator[59] ), .CK (n_0_0), .D (n_0_384));
DFF_X1 \accumulator_reg[60]  (.Q (\accumulator[60] ), .CK (n_0_0), .D (n_0_385));
DFF_X1 \accumulator_reg[61]  (.Q (\accumulator[61] ), .CK (n_0_0), .D (n_0_386));
DFF_X1 \accumulator_reg[62]  (.Q (\accumulator[62] ), .CK (n_0_0), .D (n_0_387));
DFF_X1 \accumulator_reg[63]  (.Q (\accumulator[63] ), .CK (n_0_0), .D (n_0_388));
CLKGATETST_X1 clk_gate_accumulator_reg (.GCK (n_0_0), .CK (clk), .E (n_0_389), .SE (1'b0 ));
DFF_X1 \outmultiplicand_reg_reg[0]  (.Q (\outmultiplicand_reg[0] ), .CK (n_0_1), .D (n_0_421));
DFF_X1 \outmultiplicand_reg_reg[1]  (.Q (\outmultiplicand_reg[1] ), .CK (n_0_1), .D (n_0_422));
DFF_X1 \outmultiplicand_reg_reg[2]  (.Q (\outmultiplicand_reg[2] ), .CK (n_0_1), .D (n_0_423));
DFF_X1 \outmultiplicand_reg_reg[3]  (.Q (\outmultiplicand_reg[3] ), .CK (n_0_1), .D (n_0_424));
DFF_X1 \outmultiplicand_reg_reg[4]  (.Q (\outmultiplicand_reg[4] ), .CK (n_0_1), .D (n_0_425));
DFF_X1 \outmultiplicand_reg_reg[5]  (.Q (\outmultiplicand_reg[5] ), .CK (n_0_1), .D (n_0_426));
DFF_X1 \outmultiplicand_reg_reg[6]  (.Q (\outmultiplicand_reg[6] ), .CK (n_0_1), .D (n_0_427));
DFF_X1 \outmultiplicand_reg_reg[7]  (.Q (\outmultiplicand_reg[7] ), .CK (n_0_1), .D (n_0_428));
DFF_X1 \outmultiplicand_reg_reg[8]  (.Q (\outmultiplicand_reg[8] ), .CK (n_0_1), .D (n_0_429));
DFF_X1 \outmultiplicand_reg_reg[9]  (.Q (\outmultiplicand_reg[9] ), .CK (n_0_1), .D (n_0_430));
DFF_X1 \outmultiplicand_reg_reg[10]  (.Q (\outmultiplicand_reg[10] ), .CK (n_0_1), .D (n_0_431));
DFF_X1 \outmultiplicand_reg_reg[11]  (.Q (\outmultiplicand_reg[11] ), .CK (n_0_1), .D (n_0_432));
DFF_X1 \outmultiplicand_reg_reg[12]  (.Q (\outmultiplicand_reg[12] ), .CK (n_0_1), .D (n_0_433));
DFF_X1 \outmultiplicand_reg_reg[13]  (.Q (\outmultiplicand_reg[13] ), .CK (n_0_1), .D (n_0_434));
DFF_X1 \outmultiplicand_reg_reg[14]  (.Q (\outmultiplicand_reg[14] ), .CK (n_0_1), .D (n_0_435));
DFF_X1 \outmultiplicand_reg_reg[15]  (.Q (\outmultiplicand_reg[15] ), .CK (n_0_1), .D (n_0_436));
DFF_X1 \outmultiplicand_reg_reg[16]  (.Q (\outmultiplicand_reg[16] ), .CK (n_0_1), .D (n_0_437));
DFF_X1 \outmultiplicand_reg_reg[17]  (.Q (\outmultiplicand_reg[17] ), .CK (n_0_1), .D (n_0_438));
DFF_X1 \outmultiplicand_reg_reg[18]  (.Q (\outmultiplicand_reg[18] ), .CK (n_0_1), .D (n_0_439));
DFF_X1 \outmultiplicand_reg_reg[19]  (.Q (\outmultiplicand_reg[19] ), .CK (n_0_1), .D (n_0_440));
DFF_X1 \outmultiplicand_reg_reg[20]  (.Q (\outmultiplicand_reg[20] ), .CK (n_0_1), .D (n_0_441));
DFF_X1 \outmultiplicand_reg_reg[21]  (.Q (\outmultiplicand_reg[21] ), .CK (n_0_1), .D (n_0_442));
DFF_X1 \outmultiplicand_reg_reg[22]  (.Q (\outmultiplicand_reg[22] ), .CK (n_0_1), .D (n_0_443));
DFF_X1 \outmultiplicand_reg_reg[23]  (.Q (\outmultiplicand_reg[23] ), .CK (n_0_1), .D (n_0_444));
DFF_X1 \outmultiplicand_reg_reg[24]  (.Q (\outmultiplicand_reg[24] ), .CK (n_0_1), .D (n_0_445));
DFF_X1 \outmultiplicand_reg_reg[25]  (.Q (\outmultiplicand_reg[25] ), .CK (n_0_1), .D (n_0_446));
DFF_X1 \outmultiplicand_reg_reg[26]  (.Q (\outmultiplicand_reg[26] ), .CK (n_0_1), .D (n_0_447));
DFF_X1 \outmultiplicand_reg_reg[27]  (.Q (\outmultiplicand_reg[27] ), .CK (n_0_1), .D (n_0_448));
DFF_X1 \outmultiplicand_reg_reg[28]  (.Q (\outmultiplicand_reg[28] ), .CK (n_0_1), .D (n_0_449));
DFF_X1 \outmultiplicand_reg_reg[29]  (.Q (\outmultiplicand_reg[29] ), .CK (n_0_1), .D (n_0_450));
DFF_X1 \outmultiplicand_reg_reg[30]  (.Q (\outmultiplicand_reg[30] ), .CK (n_0_1), .D (n_0_451));
DFF_X1 \outmultiplicand_reg_reg[31]  (.Q (\outmultiplicand_reg[31] ), .CK (n_0_1), .D (n_0_452));
OAI22_X1 i_0_2_667 (.ZN (n_0_323), .A1 (n_0_2_471), .A2 (n_0_2_472), .B1 (n_0_2_469), .B2 (spw__n324));
OAI21_X1 i_0_2_666 (.ZN (n_0_2_472), .A (spw__n324), .B1 (n_0_2_457), .B2 (n_0_2_150));
OAI221_X1 i_0_2_665 (.ZN (n_0_2_471), .A (n_0_2_470), .B1 (n_0_2_153), .B2 (n_0_2_449)
    , .C1 (n_0_2_155), .C2 (n_0_2_463));
OAI221_X1 i_0_2_664 (.ZN (n_0_2_470), .A (n_0_2_11), .B1 (n_0_2_341), .B2 (n_0_2_418)
    , .C1 (n_0_2_339), .C2 (n_0_2_444));
OAI22_X1 i_0_2_663 (.ZN (n_0_322), .A1 (n_0_2_464), .A2 (spw__n324), .B1 (sps__n10), .B2 (n_0_2_469));
OAI211_X1 i_0_2_662 (.ZN (n_0_2_469), .A (n_0_2_465), .B (n_0_2_468), .C1 (n_0_2_153), .C2 (n_0_2_445));
AOI22_X1 i_0_2_661 (.ZN (n_0_2_468), .A1 (n_0_2_454), .A2 (n_0_2_466), .B1 (n_0_2_467), .B2 (n_0_2_192));
INV_X1 i_0_2_660 (.ZN (n_0_2_467), .A (n_0_2_461));
INV_X1 i_0_2_659 (.ZN (n_0_2_466), .A (n_0_2_150));
OAI221_X1 i_0_2_658 (.ZN (n_0_2_465), .A (n_0_2_11), .B1 (n_0_2_332), .B2 (n_0_2_444)
    , .C1 (n_0_2_334), .C2 (n_0_2_418));
OAI22_X1 i_0_2_657 (.ZN (n_0_321), .A1 (n_0_2_462), .A2 (spw__n324), .B1 (n_0_2_464), .B2 (sps__n10));
OAI222_X1 i_0_2_656 (.ZN (n_0_2_464), .A1 (n_0_2_459), .A2 (sps__n1), .B1 (n_0_2_463)
    , .B2 (n_0_2_12), .C1 (n_0_2_449), .C2 (n_0_2_150));
OAI22_X1 i_0_2_655 (.ZN (n_0_2_463), .A1 (n_0_2_325), .A2 (n_0_2_444), .B1 (n_0_2_327), .B2 (n_0_2_418));
OAI22_X1 i_0_2_654 (.ZN (n_0_320), .A1 (n_0_2_462), .A2 (sps__n10), .B1 (spw__n326), .B2 (n_0_2_460));
OAI222_X1 i_0_2_653 (.ZN (n_0_2_462), .A1 (n_0_2_455), .A2 (sps__n1), .B1 (n_0_2_445)
    , .B2 (n_0_2_150), .C1 (n_0_2_461), .C2 (n_0_2_12));
OAI22_X1 i_0_2_652 (.ZN (n_0_2_461), .A1 (n_0_2_318), .A2 (n_0_2_444), .B1 (n_0_2_320), .B2 (n_0_2_418));
OAI22_X1 i_0_2_651 (.ZN (n_0_319), .A1 (n_0_2_456), .A2 (spw__n326), .B1 (n_0_2_460), .B2 (sps__n10));
AOI22_X1 i_0_2_650 (.ZN (n_0_2_460), .A1 (spw__n155), .A2 (n_0_2_459), .B1 (n_0_2_451), .B2 (spw__n312));
AOI22_X1 i_0_2_649 (.ZN (n_0_2_459), .A1 (n_0_2_441), .A2 (spw__n337), .B1 (n_0_2_458), .B2 (n_0_2_154));
INV_X1 i_0_2_648 (.ZN (n_0_2_458), .A (n_0_2_457));
OAI22_X1 i_0_2_647 (.ZN (n_0_2_457), .A1 (n_0_2_313), .A2 (n_0_2_418), .B1 (n_0_2_311), .B2 (n_0_2_444));
OAI22_X1 i_0_2_646 (.ZN (n_0_318), .A1 (n_0_2_452), .A2 (spw__n326), .B1 (n_0_2_456), .B2 (sps__n10));
AOI22_X1 i_0_2_645 (.ZN (n_0_2_456), .A1 (spw__n155), .A2 (n_0_2_455), .B1 (n_0_2_447), .B2 (spw__n312));
AOI22_X1 i_0_2_644 (.ZN (n_0_2_455), .A1 (n_0_2_438), .A2 (spw__n337), .B1 (n_0_2_454), .B2 (n_0_2_154));
AOI22_X1 i_0_2_643 (.ZN (n_0_2_454), .A1 (n_0_2_307), .A2 (n_0_2_419), .B1 (n_0_2_305), .B2 (n_0_2_453));
INV_X1 i_0_2_642 (.ZN (n_0_2_453), .A (n_0_2_444));
OAI22_X1 i_0_2_641 (.ZN (n_0_317), .A1 (n_0_2_448), .A2 (spw__n326), .B1 (n_0_2_452), .B2 (sps__n10));
AOI22_X1 i_0_2_640 (.ZN (n_0_2_452), .A1 (n_0_2_442), .A2 (spw__n312), .B1 (n_0_2_451), .B2 (spw__n155));
OAI22_X1 i_0_2_639 (.ZN (n_0_2_451), .A1 (n_0_2_435), .A2 (n_0_2_154), .B1 (n_0_2_450), .B2 (spw__n337));
INV_X1 i_0_2_638 (.ZN (n_0_2_450), .A (n_0_2_449));
OAI22_X1 i_0_2_637 (.ZN (n_0_2_449), .A1 (n_0_2_300), .A2 (n_0_2_418), .B1 (n_0_2_298), .B2 (n_0_2_444));
OAI22_X1 i_0_2_636 (.ZN (n_0_316), .A1 (n_0_2_443), .A2 (spw__n326), .B1 (n_0_2_448), .B2 (sps__n10));
AOI22_X1 i_0_2_635 (.ZN (n_0_2_448), .A1 (n_0_2_439), .A2 (spw__n312), .B1 (n_0_2_447), .B2 (spw__n155));
OAI22_X1 i_0_2_634 (.ZN (n_0_2_447), .A1 (n_0_2_432), .A2 (n_0_2_154), .B1 (n_0_2_446), .B2 (spw__n337));
INV_X1 i_0_2_633 (.ZN (n_0_2_446), .A (n_0_2_445));
OAI22_X1 i_0_2_632 (.ZN (n_0_2_445), .A1 (n_0_2_290), .A2 (n_0_2_444), .B1 (n_0_2_293), .B2 (n_0_2_418));
NAND2_X1 i_0_2_631 (.ZN (n_0_2_444), .A1 (\counter[5] ), .A2 (spc__n22));
OAI22_X1 i_0_2_630 (.ZN (n_0_315), .A1 (n_0_2_440), .A2 (spw__n326), .B1 (n_0_2_443), .B2 (sps__n10));
AOI22_X1 i_0_2_629 (.ZN (n_0_2_443), .A1 (n_0_2_436), .A2 (spw__n312), .B1 (n_0_2_442), .B2 (spw__n155));
OAI22_X1 i_0_2_628 (.ZN (n_0_2_442), .A1 (n_0_2_429), .A2 (n_0_2_154), .B1 (n_0_2_441), .B2 (spw__n337));
AOI22_X1 i_0_2_627 (.ZN (n_0_2_441), .A1 (n_0_2_414), .A2 (spc__n22), .B1 (n_0_2_340), .B2 (n_0_2_419));
OAI22_X1 i_0_2_626 (.ZN (n_0_314), .A1 (n_0_2_437), .A2 (spw__n326), .B1 (n_0_2_440), .B2 (sps__n10));
AOI22_X1 i_0_2_625 (.ZN (n_0_2_440), .A1 (n_0_2_433), .A2 (spw__n312), .B1 (n_0_2_439), .B2 (spw__n156));
OAI22_X1 i_0_2_624 (.ZN (n_0_2_439), .A1 (n_0_2_426), .A2 (n_0_2_154), .B1 (n_0_2_438), .B2 (spw__n337));
AOI22_X1 i_0_2_623 (.ZN (n_0_2_438), .A1 (n_0_2_409), .A2 (spc__n22), .B1 (n_0_2_333), .B2 (n_0_2_419));
OAI22_X1 i_0_2_622 (.ZN (n_0_313), .A1 (n_0_2_434), .A2 (spw__n326), .B1 (n_0_2_437), .B2 (sps__n10));
AOI22_X1 i_0_2_621 (.ZN (n_0_2_437), .A1 (n_0_2_430), .A2 (spw__n312), .B1 (n_0_2_436), .B2 (spw__n156));
OAI22_X1 i_0_2_620 (.ZN (n_0_2_436), .A1 (n_0_2_423), .A2 (n_0_2_154), .B1 (n_0_2_435), .B2 (spw__n337));
AOI22_X1 i_0_2_619 (.ZN (n_0_2_435), .A1 (n_0_2_404), .A2 (spc__n22), .B1 (n_0_2_326), .B2 (n_0_2_419));
OAI22_X1 i_0_2_618 (.ZN (n_0_312), .A1 (n_0_2_431), .A2 (spw__n325), .B1 (n_0_2_434), .B2 (sps__n10));
AOI22_X1 i_0_2_617 (.ZN (n_0_2_434), .A1 (n_0_2_427), .A2 (spw__n312), .B1 (n_0_2_433), .B2 (spw__n156));
OAI22_X1 i_0_2_616 (.ZN (n_0_2_433), .A1 (n_0_2_420), .A2 (n_0_2_154), .B1 (n_0_2_432), .B2 (spw__n338));
AOI22_X1 i_0_2_615 (.ZN (n_0_2_432), .A1 (n_0_2_399), .A2 (spc__n22), .B1 (n_0_2_319), .B2 (n_0_2_419));
OAI22_X1 i_0_2_614 (.ZN (n_0_311), .A1 (n_0_2_428), .A2 (spw__n325), .B1 (n_0_2_431), .B2 (sps__n10));
AOI22_X1 i_0_2_613 (.ZN (n_0_2_431), .A1 (n_0_2_424), .A2 (spw__n311), .B1 (n_0_2_430), .B2 (spw__n156));
OAI22_X1 i_0_2_612 (.ZN (n_0_2_430), .A1 (n_0_2_415), .A2 (n_0_2_154), .B1 (n_0_2_429), .B2 (spw__n338));
AOI22_X1 i_0_2_611 (.ZN (n_0_2_429), .A1 (n_0_2_394), .A2 (spc__n22), .B1 (n_0_2_312), .B2 (n_0_2_419));
OAI22_X1 i_0_2_610 (.ZN (n_0_310), .A1 (n_0_2_425), .A2 (spw__n325), .B1 (n_0_2_428), .B2 (sps__n10));
AOI22_X1 i_0_2_609 (.ZN (n_0_2_428), .A1 (n_0_2_421), .A2 (spw__n311), .B1 (n_0_2_427), .B2 (spw__n156));
OAI22_X1 i_0_2_608 (.ZN (n_0_2_427), .A1 (n_0_2_410), .A2 (n_0_2_154), .B1 (n_0_2_426), .B2 (spw__n338));
AOI22_X1 i_0_2_607 (.ZN (n_0_2_426), .A1 (n_0_2_389), .A2 (spc__n22), .B1 (n_0_2_305), .B2 (n_0_2_419));
OAI22_X1 i_0_2_606 (.ZN (n_0_309), .A1 (n_0_2_422), .A2 (spw__n325), .B1 (n_0_2_425), .B2 (sps__n10));
AOI22_X1 i_0_2_605 (.ZN (n_0_2_425), .A1 (n_0_2_416), .A2 (spw__n311), .B1 (n_0_2_424), .B2 (spw__n156));
OAI22_X1 i_0_2_604 (.ZN (n_0_2_424), .A1 (n_0_2_405), .A2 (n_0_2_154), .B1 (n_0_2_423), .B2 (spw__n338));
AOI22_X1 i_0_2_603 (.ZN (n_0_2_423), .A1 (n_0_2_385), .A2 (spc__n22), .B1 (n_0_2_299), .B2 (n_0_2_419));
OAI22_X1 i_0_2_602 (.ZN (n_0_308), .A1 (n_0_2_417), .A2 (spw__n325), .B1 (n_0_2_422), .B2 (sps__n10));
AOI22_X1 i_0_2_601 (.ZN (n_0_2_422), .A1 (n_0_2_411), .A2 (spw__n311), .B1 (n_0_2_421), .B2 (spw__n156));
OAI22_X1 i_0_2_600 (.ZN (n_0_2_421), .A1 (n_0_2_400), .A2 (n_0_2_154), .B1 (n_0_2_420), .B2 (spw__n338));
AOI22_X1 i_0_2_599 (.ZN (n_0_2_420), .A1 (n_0_2_380), .A2 (spc__n22), .B1 (n_0_2_291), .B2 (n_0_2_419));
INV_X1 i_0_2_598 (.ZN (n_0_2_419), .A (n_0_2_418));
NAND2_X1 i_0_2_597 (.ZN (n_0_2_418), .A1 (spc__n19), .A2 (\counter[5] ));
OAI22_X1 i_0_2_596 (.ZN (n_0_307), .A1 (n_0_2_412), .A2 (spw__n325), .B1 (n_0_2_417), .B2 (sps__n10));
AOI22_X1 i_0_2_595 (.ZN (n_0_2_417), .A1 (n_0_2_406), .A2 (spw__n311), .B1 (n_0_2_416), .B2 (spw__n156));
OAI22_X1 i_0_2_594 (.ZN (n_0_2_416), .A1 (n_0_2_415), .A2 (spw__n338), .B1 (n_0_2_395), .B2 (n_0_2_154));
AOI22_X1 i_0_2_593 (.ZN (n_0_2_415), .A1 (n_0_2_375), .A2 (spc__n22), .B1 (n_0_2_414), .B2 (spc__n19));
OAI22_X1 i_0_2_592 (.ZN (n_0_2_414), .A1 (n_0_2_14), .A2 (n_0_2_284), .B1 (n_0_2_346), .B2 (n_0_2_413));
INV_X1 i_0_2_591 (.ZN (n_0_2_413), .A (\multiplicand1[31] ));
OAI22_X1 i_0_2_590 (.ZN (n_0_306), .A1 (n_0_2_412), .A2 (sps__n10), .B1 (n_0_2_407), .B2 (spw__n325));
AOI22_X1 i_0_2_589 (.ZN (n_0_2_412), .A1 (n_0_2_401), .A2 (spw__n310), .B1 (n_0_2_411), .B2 (spw__n156));
OAI22_X1 i_0_2_588 (.ZN (n_0_2_411), .A1 (n_0_2_410), .A2 (spw__n338), .B1 (n_0_2_390), .B2 (n_0_2_154));
AOI22_X1 i_0_2_587 (.ZN (n_0_2_410), .A1 (n_0_2_371), .A2 (spc__n22), .B1 (n_0_2_409), .B2 (spc__n19));
OAI22_X1 i_0_2_586 (.ZN (n_0_2_409), .A1 (n_0_2_14), .A2 (n_0_2_278), .B1 (n_0_2_346), .B2 (n_0_2_408));
INV_X1 i_0_2_585 (.ZN (n_0_2_408), .A (\multiplicand1[30] ));
OAI22_X1 i_0_2_584 (.ZN (n_0_305), .A1 (n_0_2_402), .A2 (spw__n325), .B1 (n_0_2_407), .B2 (sps__n10));
AOI22_X1 i_0_2_583 (.ZN (n_0_2_407), .A1 (n_0_2_406), .A2 (spw__n156), .B1 (n_0_2_396), .B2 (spw__n310));
OAI22_X1 i_0_2_582 (.ZN (n_0_2_406), .A1 (n_0_2_405), .A2 (spw__n338), .B1 (n_0_2_386), .B2 (n_0_2_154));
AOI22_X1 i_0_2_581 (.ZN (n_0_2_405), .A1 (n_0_2_367), .A2 (spc__n22), .B1 (n_0_2_404), .B2 (spc__n19));
OAI22_X1 i_0_2_580 (.ZN (n_0_2_404), .A1 (n_0_2_14), .A2 (n_0_2_272), .B1 (n_0_2_346), .B2 (n_0_2_403));
INV_X1 i_0_2_579 (.ZN (n_0_2_403), .A (\multiplicand1[29] ));
OAI22_X1 i_0_2_578 (.ZN (n_0_304), .A1 (n_0_2_402), .A2 (sps__n10), .B1 (n_0_2_397), .B2 (spw__n325));
AOI22_X1 i_0_2_577 (.ZN (n_0_2_402), .A1 (n_0_2_401), .A2 (spw__n156), .B1 (n_0_2_391), .B2 (spw__n310));
OAI22_X1 i_0_2_576 (.ZN (n_0_2_401), .A1 (n_0_2_400), .A2 (spw__n338), .B1 (n_0_2_381), .B2 (n_0_2_154));
AOI22_X1 i_0_2_575 (.ZN (n_0_2_400), .A1 (n_0_2_363), .A2 (spc__n22), .B1 (n_0_2_399), .B2 (spc__n19));
OAI22_X1 i_0_2_574 (.ZN (n_0_2_399), .A1 (n_0_2_14), .A2 (n_0_2_265), .B1 (n_0_2_346), .B2 (n_0_2_398));
INV_X1 i_0_2_573 (.ZN (n_0_2_398), .A (\multiplicand1[28] ));
OAI22_X1 i_0_2_572 (.ZN (n_0_303), .A1 (n_0_2_392), .A2 (spw__n325), .B1 (n_0_2_397), .B2 (sps__n10));
AOI22_X1 i_0_2_571 (.ZN (n_0_2_397), .A1 (n_0_2_387), .A2 (spw__n310), .B1 (n_0_2_396), .B2 (spw__n156));
OAI22_X1 i_0_2_570 (.ZN (n_0_2_396), .A1 (n_0_2_395), .A2 (spw__n338), .B1 (n_0_2_376), .B2 (n_0_2_154));
AOI22_X1 i_0_2_569 (.ZN (n_0_2_395), .A1 (n_0_2_394), .A2 (spc__n19), .B1 (n_0_2_359), .B2 (spc__n22));
OAI22_X1 i_0_2_568 (.ZN (n_0_2_394), .A1 (n_0_2_14), .A2 (n_0_2_225), .B1 (n_0_2_346), .B2 (n_0_2_393));
INV_X1 i_0_2_567 (.ZN (n_0_2_393), .A (\multiplicand1[27] ));
OAI22_X1 i_0_2_566 (.ZN (n_0_302), .A1 (n_0_2_392), .A2 (sps__n10), .B1 (n_0_2_388), .B2 (spw__n325));
AOI22_X1 i_0_2_565 (.ZN (n_0_2_392), .A1 (n_0_2_382), .A2 (spw__n310), .B1 (n_0_2_391), .B2 (spw__n156));
OAI22_X1 i_0_2_564 (.ZN (n_0_2_391), .A1 (n_0_2_390), .A2 (spw__n338), .B1 (n_0_2_372), .B2 (n_0_2_154));
AOI22_X1 i_0_2_563 (.ZN (n_0_2_390), .A1 (n_0_2_389), .A2 (spc__n19), .B1 (n_0_2_355), .B2 (spc__n22));
OAI22_X1 i_0_2_562 (.ZN (n_0_2_389), .A1 (n_0_2_14), .A2 (n_0_2_218), .B1 (n_0_2_346), .B2 (n_0_2_306));
OAI22_X1 i_0_2_561 (.ZN (n_0_301), .A1 (n_0_2_383), .A2 (spw__n325), .B1 (n_0_2_388), .B2 (sps__n10));
AOI22_X1 i_0_2_560 (.ZN (n_0_2_388), .A1 (n_0_2_387), .A2 (spw__n156), .B1 (n_0_2_377), .B2 (spw__n310));
OAI22_X1 i_0_2_559 (.ZN (n_0_2_387), .A1 (n_0_2_386), .A2 (spw__n338), .B1 (n_0_2_368), .B2 (n_0_2_154));
AOI22_X1 i_0_2_558 (.ZN (n_0_2_386), .A1 (n_0_2_385), .A2 (spc__n19), .B1 (n_0_2_351), .B2 (spc__n22));
OAI22_X1 i_0_2_557 (.ZN (n_0_2_385), .A1 (n_0_2_14), .A2 (n_0_2_249), .B1 (n_0_2_346), .B2 (n_0_2_384));
INV_X1 i_0_2_556 (.ZN (n_0_2_384), .A (\multiplicand1[25] ));
OAI22_X1 i_0_2_555 (.ZN (n_0_300), .A1 (n_0_2_383), .A2 (sps__n10), .B1 (n_0_2_378), .B2 (spw__n325));
AOI22_X1 i_0_2_554 (.ZN (n_0_2_383), .A1 (n_0_2_382), .A2 (spw__n156), .B1 (n_0_2_373), .B2 (spw__n310));
OAI22_X1 i_0_2_553 (.ZN (n_0_2_382), .A1 (n_0_2_381), .A2 (spw__n338), .B1 (n_0_2_364), .B2 (n_0_2_154));
AOI22_X1 i_0_2_552 (.ZN (n_0_2_381), .A1 (n_0_2_380), .A2 (spc__n19), .B1 (n_0_2_347), .B2 (spc__n22));
OAI22_X1 i_0_2_551 (.ZN (n_0_2_380), .A1 (n_0_2_14), .A2 (n_0_2_242), .B1 (n_0_2_346), .B2 (n_0_2_379));
INV_X1 i_0_2_550 (.ZN (n_0_2_379), .A (\multiplicand1[24] ));
OAI22_X1 i_0_2_549 (.ZN (n_0_299), .A1 (n_0_2_374), .A2 (spw__n325), .B1 (n_0_2_378), .B2 (sps__n10));
AOI22_X1 i_0_2_548 (.ZN (n_0_2_378), .A1 (n_0_2_369), .A2 (spw__n310), .B1 (n_0_2_377), .B2 (spw__n156));
OAI22_X1 i_0_2_547 (.ZN (n_0_2_377), .A1 (n_0_2_376), .A2 (spw__n338), .B1 (n_0_2_360), .B2 (n_0_2_154));
AOI22_X1 i_0_2_546 (.ZN (n_0_2_376), .A1 (n_0_2_375), .A2 (spc__n19), .B1 (n_0_2_342), .B2 (n_0_2_292));
OAI22_X1 i_0_2_545 (.ZN (n_0_2_375), .A1 (n_0_2_14), .A2 (n_0_2_204), .B1 (n_0_2_346), .B2 (n_0_2_285));
OAI22_X1 i_0_2_544 (.ZN (n_0_298), .A1 (n_0_2_374), .A2 (sps__n10), .B1 (n_0_2_370), .B2 (spw__n325));
AOI22_X1 i_0_2_543 (.ZN (n_0_2_374), .A1 (n_0_2_365), .A2 (spw__n310), .B1 (n_0_2_373), .B2 (spw__n156));
OAI22_X1 i_0_2_542 (.ZN (n_0_2_373), .A1 (n_0_2_372), .A2 (spw__n338), .B1 (n_0_2_356), .B2 (n_0_2_154));
AOI22_X1 i_0_2_541 (.ZN (n_0_2_372), .A1 (n_0_2_371), .A2 (spc__n19), .B1 (n_0_2_335), .B2 (n_0_2_292));
OAI22_X1 i_0_2_540 (.ZN (n_0_2_371), .A1 (n_0_2_14), .A2 (n_0_2_199), .B1 (n_0_2_346), .B2 (n_0_2_279));
OAI22_X1 i_0_2_539 (.ZN (n_0_297), .A1 (n_0_2_366), .A2 (spw__n325), .B1 (n_0_2_370), .B2 (sps__n10));
AOI22_X1 i_0_2_538 (.ZN (n_0_2_370), .A1 (n_0_2_369), .A2 (spw__n156), .B1 (n_0_2_361), .B2 (spw__n310));
OAI22_X1 i_0_2_537 (.ZN (n_0_2_369), .A1 (n_0_2_368), .A2 (spw__n338), .B1 (n_0_2_352), .B2 (n_0_2_154));
AOI22_X1 i_0_2_536 (.ZN (n_0_2_368), .A1 (n_0_2_367), .A2 (spc__n19), .B1 (n_0_2_328), .B2 (n_0_2_292));
OAI22_X1 i_0_2_535 (.ZN (n_0_2_367), .A1 (n_0_2_14), .A2 (n_0_2_195), .B1 (n_0_2_346), .B2 (n_0_2_273));
OAI22_X1 i_0_2_534 (.ZN (n_0_296), .A1 (n_0_2_366), .A2 (sps__n10), .B1 (n_0_2_362), .B2 (spw__n325));
AOI22_X1 i_0_2_533 (.ZN (n_0_2_366), .A1 (n_0_2_365), .A2 (spw__n156), .B1 (n_0_2_357), .B2 (spw__n310));
OAI22_X1 i_0_2_532 (.ZN (n_0_2_365), .A1 (n_0_2_364), .A2 (spw__n338), .B1 (n_0_2_348), .B2 (n_0_2_154));
AOI22_X1 i_0_2_531 (.ZN (n_0_2_364), .A1 (n_0_2_363), .A2 (spc__n19), .B1 (n_0_2_321), .B2 (n_0_2_292));
OAI22_X1 i_0_2_530 (.ZN (n_0_2_363), .A1 (n_0_2_14), .A2 (n_0_2_190), .B1 (n_0_2_346), .B2 (n_0_2_266));
OAI22_X1 i_0_2_529 (.ZN (n_0_295), .A1 (n_0_2_358), .A2 (spw__n325), .B1 (n_0_2_362), .B2 (sps__n10));
AOI22_X1 i_0_2_528 (.ZN (n_0_2_362), .A1 (n_0_2_353), .A2 (spw__n311), .B1 (n_0_2_361), .B2 (spw__n156));
OAI22_X1 i_0_2_527 (.ZN (n_0_2_361), .A1 (n_0_2_360), .A2 (spw__n338), .B1 (n_0_2_343), .B2 (n_0_2_154));
AOI22_X1 i_0_2_526 (.ZN (n_0_2_360), .A1 (n_0_2_359), .A2 (spc__n19), .B1 (n_0_2_314), .B2 (n_0_2_292));
OAI22_X1 i_0_2_525 (.ZN (n_0_2_359), .A1 (n_0_2_346), .A2 (n_0_2_260), .B1 (n_0_2_14), .B2 (n_0_2_203));
OAI22_X1 i_0_2_524 (.ZN (n_0_294), .A1 (n_0_2_358), .A2 (sps__n10), .B1 (n_0_2_354), .B2 (spw__n325));
AOI22_X1 i_0_2_523 (.ZN (n_0_2_358), .A1 (n_0_2_349), .A2 (spw__n311), .B1 (n_0_2_357), .B2 (spw__n156));
OAI22_X1 i_0_2_522 (.ZN (n_0_2_357), .A1 (n_0_2_356), .A2 (spw__n338), .B1 (n_0_2_336), .B2 (n_0_2_154));
AOI22_X1 i_0_2_521 (.ZN (n_0_2_356), .A1 (n_0_2_355), .A2 (spc__n19), .B1 (n_0_2_307), .B2 (n_0_2_292));
OAI22_X1 i_0_2_520 (.ZN (n_0_2_355), .A1 (n_0_2_346), .A2 (n_0_2_255), .B1 (n_0_2_14), .B2 (n_0_2_198));
OAI22_X1 i_0_2_519 (.ZN (n_0_293), .A1 (n_0_2_350), .A2 (spw__n325), .B1 (n_0_2_354), .B2 (sps__n10));
AOI22_X1 i_0_2_518 (.ZN (n_0_2_354), .A1 (n_0_2_353), .A2 (spw__n156), .B1 (n_0_2_344), .B2 (spw__n312));
OAI22_X1 i_0_2_517 (.ZN (n_0_2_353), .A1 (n_0_2_352), .A2 (spw__n338), .B1 (n_0_2_329), .B2 (n_0_2_154));
AOI22_X1 i_0_2_516 (.ZN (n_0_2_352), .A1 (n_0_2_351), .A2 (spc__n19), .B1 (n_0_2_301), .B2 (n_0_2_292));
OAI22_X1 i_0_2_515 (.ZN (n_0_2_351), .A1 (n_0_2_14), .A2 (n_0_2_185), .B1 (n_0_2_346), .B2 (n_0_2_250));
OAI22_X1 i_0_2_514 (.ZN (n_0_292), .A1 (n_0_2_350), .A2 (sps__n10), .B1 (n_0_2_345), .B2 (spw__n325));
AOI22_X1 i_0_2_513 (.ZN (n_0_2_350), .A1 (n_0_2_349), .A2 (spw__n156), .B1 (n_0_2_337), .B2 (spw__n312));
OAI22_X1 i_0_2_512 (.ZN (n_0_2_349), .A1 (n_0_2_348), .A2 (spw__n338), .B1 (n_0_2_322), .B2 (n_0_2_154));
AOI22_X1 i_0_2_511 (.ZN (n_0_2_348), .A1 (n_0_2_347), .A2 (spc__n19), .B1 (n_0_2_294), .B2 (n_0_2_292));
OAI22_X1 i_0_2_510 (.ZN (n_0_2_347), .A1 (n_0_2_14), .A2 (n_0_2_183), .B1 (n_0_2_346), .B2 (n_0_2_243));
NAND2_X1 i_0_2_509 (.ZN (n_0_2_346), .A1 (n_0_2_10), .A2 (spc__n16));
OAI22_X1 i_0_2_508 (.ZN (n_0_291), .A1 (n_0_2_338), .A2 (spw__n324), .B1 (n_0_2_345), .B2 (sps__n10));
AOI22_X1 i_0_2_507 (.ZN (n_0_2_345), .A1 (n_0_2_330), .A2 (spw__n309), .B1 (n_0_2_344), .B2 (spw__n155));
OAI22_X1 i_0_2_506 (.ZN (n_0_2_344), .A1 (n_0_2_315), .A2 (n_0_2_154), .B1 (n_0_2_343), .B2 (spw__n337));
AOI22_X1 i_0_2_505 (.ZN (n_0_2_343), .A1 (n_0_2_340), .A2 (n_0_2_292), .B1 (n_0_2_342), .B2 (n_0_2_180));
INV_X1 i_0_2_504 (.ZN (n_0_2_342), .A (n_0_2_341));
OAI22_X1 i_0_2_503 (.ZN (n_0_2_341), .A1 (n_0_2_13), .A2 (\multiplicand1[15] ), .B1 (spc__n16), .B2 (\multiplicand1[31] ));
INV_X1 i_0_2_502 (.ZN (n_0_2_340), .A (n_0_2_339));
OAI22_X1 i_0_2_501 (.ZN (n_0_2_339), .A1 (n_0_2_13), .A2 (\multiplicand1[7] ), .B1 (spc__n16), .B2 (\multiplicand1[23] ));
OAI22_X1 i_0_2_500 (.ZN (n_0_290), .A1 (n_0_2_331), .A2 (spw__n324), .B1 (sps__n10), .B2 (n_0_2_338));
AOI22_X1 i_0_2_499 (.ZN (n_0_2_338), .A1 (n_0_2_323), .A2 (spw__n309), .B1 (n_0_2_337), .B2 (spw__n155));
OAI22_X1 i_0_2_498 (.ZN (n_0_2_337), .A1 (n_0_2_308), .A2 (n_0_2_154), .B1 (n_0_2_336), .B2 (spw__n337));
AOI22_X1 i_0_2_497 (.ZN (n_0_2_336), .A1 (n_0_2_333), .A2 (n_0_2_292), .B1 (n_0_2_335), .B2 (n_0_2_180));
INV_X1 i_0_2_496 (.ZN (n_0_2_335), .A (n_0_2_334));
OAI22_X1 i_0_2_495 (.ZN (n_0_2_334), .A1 (n_0_2_13), .A2 (\multiplicand1[14] ), .B1 (spc__n16), .B2 (\multiplicand1[30] ));
INV_X1 i_0_2_494 (.ZN (n_0_2_333), .A (n_0_2_332));
OAI22_X1 i_0_2_493 (.ZN (n_0_2_332), .A1 (n_0_2_13), .A2 (\multiplicand1[6] ), .B1 (spc__n16), .B2 (\multiplicand1[22] ));
OAI22_X1 i_0_2_492 (.ZN (n_0_289), .A1 (n_0_2_324), .A2 (spw__n324), .B1 (n_0_2_331), .B2 (sps__n10));
AOI22_X1 i_0_2_491 (.ZN (n_0_2_331), .A1 (n_0_2_316), .A2 (spw__n309), .B1 (spw__n155), .B2 (n_0_2_330));
OAI22_X1 i_0_2_490 (.ZN (n_0_2_330), .A1 (n_0_2_302), .A2 (n_0_2_154), .B1 (n_0_2_329), .B2 (spw__n337));
AOI22_X1 i_0_2_489 (.ZN (n_0_2_329), .A1 (n_0_2_326), .A2 (n_0_2_292), .B1 (n_0_2_328), .B2 (n_0_2_180));
INV_X1 i_0_2_488 (.ZN (n_0_2_328), .A (n_0_2_327));
OAI22_X1 i_0_2_487 (.ZN (n_0_2_327), .A1 (n_0_2_13), .A2 (\multiplicand1[13] ), .B1 (spc__n16), .B2 (\multiplicand1[29] ));
INV_X1 i_0_2_486 (.ZN (n_0_2_326), .A (n_0_2_325));
OAI22_X1 i_0_2_485 (.ZN (n_0_2_325), .A1 (n_0_2_13), .A2 (\multiplicand1[5] ), .B1 (spc__n16), .B2 (\multiplicand1[21] ));
OAI22_X1 i_0_2_484 (.ZN (n_0_288), .A1 (n_0_2_317), .A2 (spw__n324), .B1 (n_0_2_324), .B2 (sps__n10));
AOI22_X1 i_0_2_483 (.ZN (n_0_2_324), .A1 (n_0_2_309), .A2 (sps__n7), .B1 (sps__n1), .B2 (n_0_2_323));
OAI22_X1 i_0_2_482 (.ZN (n_0_2_323), .A1 (n_0_2_295), .A2 (n_0_2_154), .B1 (n_0_2_322), .B2 (spw__n337));
AOI22_X1 i_0_2_481 (.ZN (n_0_2_322), .A1 (n_0_2_319), .A2 (n_0_2_292), .B1 (n_0_2_321), .B2 (n_0_2_180));
INV_X1 i_0_2_480 (.ZN (n_0_2_321), .A (n_0_2_320));
OAI22_X1 i_0_2_479 (.ZN (n_0_2_320), .A1 (n_0_2_13), .A2 (\multiplicand1[12] ), .B1 (spc__n16), .B2 (\multiplicand1[28] ));
INV_X1 i_0_2_478 (.ZN (n_0_2_319), .A (n_0_2_318));
OAI22_X1 i_0_2_477 (.ZN (n_0_2_318), .A1 (n_0_2_13), .A2 (\multiplicand1[4] ), .B1 (spc__n16), .B2 (\multiplicand1[20] ));
OAI22_X1 i_0_2_476 (.ZN (n_0_287), .A1 (n_0_2_310), .A2 (n_0_2_148), .B1 (n_0_2_317), .B2 (sps__n10));
AOI22_X1 i_0_2_475 (.ZN (n_0_2_317), .A1 (n_0_2_303), .A2 (sps__n7), .B1 (n_0_2_316), .B2 (sps__n1));
OAI22_X1 i_0_2_474 (.ZN (n_0_2_316), .A1 (n_0_2_287), .A2 (n_0_2_269), .B1 (sps__n4), .B2 (n_0_2_315));
AOI22_X1 i_0_2_473 (.ZN (n_0_2_315), .A1 (n_0_2_312), .A2 (n_0_2_292), .B1 (n_0_2_314), .B2 (n_0_2_180));
INV_X1 i_0_2_472 (.ZN (n_0_2_314), .A (n_0_2_313));
OAI22_X1 i_0_2_471 (.ZN (n_0_2_313), .A1 (n_0_2_13), .A2 (\multiplicand1[11] ), .B1 (spc__n16), .B2 (\multiplicand1[27] ));
INV_X1 i_0_2_470 (.ZN (n_0_2_312), .A (n_0_2_311));
OAI22_X1 i_0_2_469 (.ZN (n_0_2_311), .A1 (n_0_2_13), .A2 (\multiplicand1[3] ), .B1 (spc__n16), .B2 (\multiplicand1[19] ));
OAI22_X1 i_0_2_468 (.ZN (n_0_286), .A1 (n_0_2_304), .A2 (n_0_2_148), .B1 (n_0_2_310), .B2 (sps__n10));
AOI22_X1 i_0_2_467 (.ZN (n_0_2_310), .A1 (n_0_2_296), .A2 (sps__n7), .B1 (n_0_2_309), .B2 (sps__n1));
OAI22_X1 i_0_2_466 (.ZN (n_0_2_309), .A1 (n_0_2_281), .A2 (n_0_2_269), .B1 (sps__n4), .B2 (n_0_2_308));
AOI22_X1 i_0_2_465 (.ZN (n_0_2_308), .A1 (n_0_2_305), .A2 (n_0_2_292), .B1 (n_0_2_307), .B2 (n_0_2_180));
AOI22_X1 i_0_2_464 (.ZN (n_0_2_307), .A1 (n_0_2_13), .A2 (n_0_2_306), .B1 (n_0_2_218), .B2 (spc__n16));
INV_X1 i_0_2_463 (.ZN (n_0_2_306), .A (\multiplicand1[26] ));
AOI22_X1 i_0_2_462 (.ZN (n_0_2_305), .A1 (n_0_2_13), .A2 (n_0_2_255), .B1 (n_0_2_198), .B2 (spc__n16));
OAI22_X1 i_0_2_461 (.ZN (n_0_285), .A1 (n_0_2_297), .A2 (n_0_2_148), .B1 (n_0_2_304), .B2 (sps__n10));
AOI22_X1 i_0_2_460 (.ZN (n_0_2_304), .A1 (n_0_2_288), .A2 (sps__n7), .B1 (n_0_2_303), .B2 (sps__n1));
OAI22_X1 i_0_2_459 (.ZN (n_0_2_303), .A1 (n_0_2_275), .A2 (n_0_2_269), .B1 (sps__n4), .B2 (n_0_2_302));
AOI22_X1 i_0_2_458 (.ZN (n_0_2_302), .A1 (n_0_2_299), .A2 (n_0_2_292), .B1 (n_0_2_301), .B2 (n_0_2_180));
INV_X1 i_0_2_457 (.ZN (n_0_2_301), .A (n_0_2_300));
OAI22_X1 i_0_2_456 (.ZN (n_0_2_300), .A1 (n_0_2_13), .A2 (\multiplicand1[9] ), .B1 (spc__n16), .B2 (\multiplicand1[25] ));
INV_X1 i_0_2_455 (.ZN (n_0_2_299), .A (n_0_2_298));
OAI22_X1 i_0_2_454 (.ZN (n_0_2_298), .A1 (n_0_2_13), .A2 (\multiplicand1[1] ), .B1 (spc__n16), .B2 (\multiplicand1[17] ));
OAI22_X1 i_0_2_453 (.ZN (n_0_284), .A1 (n_0_2_289), .A2 (n_0_2_148), .B1 (n_0_2_297), .B2 (sps__n10));
AOI22_X1 i_0_2_452 (.ZN (n_0_2_297), .A1 (n_0_2_282), .A2 (sps__n7), .B1 (n_0_2_296), .B2 (sps__n1));
OAI22_X1 i_0_2_451 (.ZN (n_0_2_296), .A1 (n_0_2_268), .A2 (n_0_2_269), .B1 (sps__n4), .B2 (n_0_2_295));
AOI22_X1 i_0_2_450 (.ZN (n_0_2_295), .A1 (n_0_2_291), .A2 (n_0_2_292), .B1 (n_0_2_294), .B2 (n_0_2_180));
INV_X1 i_0_2_449 (.ZN (n_0_2_294), .A (n_0_2_293));
OAI22_X1 i_0_2_448 (.ZN (n_0_2_293), .A1 (n_0_2_13), .A2 (\multiplicand1[8] ), .B1 (spc__n16), .B2 (\multiplicand1[24] ));
INV_X1 i_0_2_447 (.ZN (n_0_2_292), .A (n_0_2_219));
INV_X1 i_0_2_446 (.ZN (n_0_2_291), .A (n_0_2_290));
OAI22_X1 i_0_2_445 (.ZN (n_0_2_290), .A1 (n_0_2_13), .A2 (\multiplicand1[0] ), .B1 (spc__n16), .B2 (\multiplicand1[16] ));
OAI22_X1 i_0_2_444 (.ZN (n_0_283), .A1 (n_0_2_283), .A2 (n_0_2_148), .B1 (n_0_2_289), .B2 (sps__n10));
AOI22_X1 i_0_2_443 (.ZN (n_0_2_289), .A1 (n_0_2_276), .A2 (sps__n7), .B1 (n_0_2_288), .B2 (sps__n1));
OAI22_X1 i_0_2_442 (.ZN (n_0_2_288), .A1 (n_0_2_287), .A2 (n_0_2_246), .B1 (n_0_2_262), .B2 (n_0_2_269));
AOI21_X1 i_0_2_441 (.ZN (n_0_2_287), .A (n_0_2_286), .B1 (\multiplicand1[7] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_440 (.ZN (n_0_2_286), .A (spc__n16), .B1 (n_0_2_284), .B2 (spc__n22)
    , .C1 (n_0_2_285), .C2 (spc__n19));
INV_X1 i_0_2_439 (.ZN (n_0_2_285), .A (\multiplicand1[23] ));
INV_X1 i_0_2_438 (.ZN (n_0_2_284), .A (\multiplicand1[15] ));
OAI22_X1 i_0_2_437 (.ZN (n_0_282), .A1 (n_0_2_283), .A2 (sps__n10), .B1 (n_0_2_277), .B2 (n_0_2_148));
AOI22_X1 i_0_2_436 (.ZN (n_0_2_283), .A1 (n_0_2_270), .A2 (sps__n7), .B1 (n_0_2_282), .B2 (sps__n1));
OAI22_X1 i_0_2_435 (.ZN (n_0_2_282), .A1 (n_0_2_281), .A2 (n_0_2_246), .B1 (n_0_2_257), .B2 (n_0_2_269));
AOI21_X1 i_0_2_434 (.ZN (n_0_2_281), .A (n_0_2_280), .B1 (\multiplicand1[6] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_433 (.ZN (n_0_2_280), .A (spc__n16), .B1 (n_0_2_278), .B2 (spc__n22)
    , .C1 (n_0_2_279), .C2 (spc__n19));
INV_X1 i_0_2_432 (.ZN (n_0_2_279), .A (\multiplicand1[22] ));
INV_X1 i_0_2_431 (.ZN (n_0_2_278), .A (\multiplicand1[14] ));
OAI22_X1 i_0_2_430 (.ZN (n_0_281), .A1 (n_0_2_271), .A2 (n_0_2_148), .B1 (n_0_2_277), .B2 (sps__n10));
AOI22_X1 i_0_2_429 (.ZN (n_0_2_277), .A1 (n_0_2_276), .A2 (sps__n1), .B1 (n_0_2_263), .B2 (sps__n7));
OAI22_X1 i_0_2_428 (.ZN (n_0_2_276), .A1 (n_0_2_275), .A2 (n_0_2_246), .B1 (n_0_2_252), .B2 (n_0_2_269));
AOI21_X1 i_0_2_427 (.ZN (n_0_2_275), .A (n_0_2_274), .B1 (\multiplicand1[5] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_426 (.ZN (n_0_2_274), .A (spc__n16), .B1 (n_0_2_272), .B2 (spc__n22)
    , .C1 (n_0_2_273), .C2 (spc__n19));
INV_X1 i_0_2_425 (.ZN (n_0_2_273), .A (\multiplicand1[21] ));
INV_X1 i_0_2_424 (.ZN (n_0_2_272), .A (\multiplicand1[13] ));
OAI22_X1 i_0_2_423 (.ZN (n_0_280), .A1 (n_0_2_271), .A2 (sps__n10), .B1 (n_0_2_264), .B2 (n_0_2_148));
AOI22_X1 i_0_2_422 (.ZN (n_0_2_271), .A1 (n_0_2_270), .A2 (sps__n1), .B1 (n_0_2_258), .B2 (sps__n7));
OAI22_X1 i_0_2_421 (.ZN (n_0_2_270), .A1 (n_0_2_268), .A2 (n_0_2_246), .B1 (n_0_2_245), .B2 (n_0_2_269));
NAND2_X1 i_0_2_420 (.ZN (n_0_2_269), .A1 (n_0_2_10), .A2 (sps__n4));
AOI21_X1 i_0_2_419 (.ZN (n_0_2_268), .A (n_0_2_267), .B1 (\multiplicand1[4] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_418 (.ZN (n_0_2_267), .A (spc__n16), .B1 (n_0_2_265), .B2 (spc__n22)
    , .C1 (n_0_2_266), .C2 (spc__n19));
INV_X1 i_0_2_417 (.ZN (n_0_2_266), .A (\multiplicand1[20] ));
INV_X1 i_0_2_416 (.ZN (n_0_2_265), .A (\multiplicand1[12] ));
OAI22_X1 i_0_2_415 (.ZN (n_0_279), .A1 (n_0_2_259), .A2 (n_0_2_148), .B1 (n_0_2_264), .B2 (sps__n10));
AOI22_X1 i_0_2_414 (.ZN (n_0_2_264), .A1 (n_0_2_253), .A2 (sps__n7), .B1 (n_0_2_263), .B2 (sps__n1));
OAI22_X1 i_0_2_413 (.ZN (n_0_2_263), .A1 (n_0_2_262), .A2 (n_0_2_246), .B1 (n_0_2_239), .B2 (n_0_2_154));
AOI21_X1 i_0_2_412 (.ZN (n_0_2_262), .A (n_0_2_261), .B1 (\multiplicand1[3] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_411 (.ZN (n_0_2_261), .A (spc__n16), .B1 (n_0_2_225), .B2 (spc__n22)
    , .C1 (n_0_2_260), .C2 (spc__n19));
INV_X1 i_0_2_410 (.ZN (n_0_2_260), .A (\multiplicand1[19] ));
OAI22_X1 i_0_2_409 (.ZN (n_0_278), .A1 (n_0_2_254), .A2 (n_0_2_148), .B1 (n_0_2_259), .B2 (sps__n10));
AOI22_X1 i_0_2_408 (.ZN (n_0_2_259), .A1 (n_0_2_247), .A2 (sps__n7), .B1 (n_0_2_258), .B2 (sps__n1));
OAI22_X1 i_0_2_407 (.ZN (n_0_2_258), .A1 (n_0_2_257), .A2 (n_0_2_246), .B1 (n_0_2_236), .B2 (n_0_2_154));
AOI21_X1 i_0_2_406 (.ZN (n_0_2_257), .A (n_0_2_256), .B1 (\multiplicand1[2] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_405 (.ZN (n_0_2_256), .A (spc__n16), .B1 (n_0_2_218), .B2 (spc__n22)
    , .C1 (n_0_2_255), .C2 (spc__n19));
INV_X1 i_0_2_404 (.ZN (n_0_2_255), .A (\multiplicand1[18] ));
OAI22_X1 i_0_2_403 (.ZN (n_0_277), .A1 (n_0_2_254), .A2 (sps__n10), .B1 (n_0_2_248), .B2 (n_0_2_148));
AOI22_X1 i_0_2_402 (.ZN (n_0_2_254), .A1 (n_0_2_240), .A2 (sps__n7), .B1 (n_0_2_253), .B2 (sps__n1));
OAI22_X1 i_0_2_401 (.ZN (n_0_2_253), .A1 (n_0_2_252), .A2 (n_0_2_246), .B1 (n_0_2_233), .B2 (n_0_2_154));
AOI21_X1 i_0_2_400 (.ZN (n_0_2_252), .A (n_0_2_251), .B1 (\multiplicand1[1] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_399 (.ZN (n_0_2_251), .A (spc__n16), .B1 (n_0_2_249), .B2 (spc__n22)
    , .C1 (n_0_2_250), .C2 (spc__n19));
INV_X1 i_0_2_398 (.ZN (n_0_2_250), .A (\multiplicand1[17] ));
INV_X1 i_0_2_397 (.ZN (n_0_2_249), .A (\multiplicand1[9] ));
OAI22_X1 i_0_2_396 (.ZN (n_0_276), .A1 (n_0_2_248), .A2 (sps__n10), .B1 (n_0_2_241), .B2 (n_0_2_148));
AOI22_X1 i_0_2_395 (.ZN (n_0_2_248), .A1 (n_0_2_237), .A2 (sps__n7), .B1 (n_0_2_247), .B2 (sps__n1));
OAI22_X1 i_0_2_394 (.ZN (n_0_2_247), .A1 (n_0_2_245), .A2 (n_0_2_246), .B1 (n_0_2_230), .B2 (n_0_2_154));
NAND2_X1 i_0_2_393 (.ZN (n_0_2_246), .A1 (n_0_2_10), .A2 (n_0_2_154));
AOI21_X1 i_0_2_392 (.ZN (n_0_2_245), .A (n_0_2_244), .B1 (\multiplicand1[0] ), .B2 (n_0_2_161));
AOI221_X1 i_0_2_391 (.ZN (n_0_2_244), .A (spc__n16), .B1 (n_0_2_242), .B2 (spc__n22)
    , .C1 (n_0_2_243), .C2 (spc__n19));
INV_X1 i_0_2_390 (.ZN (n_0_2_243), .A (\multiplicand1[16] ));
INV_X1 i_0_2_389 (.ZN (n_0_2_242), .A (\multiplicand1[8] ));
OAI22_X1 i_0_2_388 (.ZN (n_0_275), .A1 (n_0_2_241), .A2 (sps__n10), .B1 (n_0_2_238), .B2 (n_0_2_148));
AOI22_X1 i_0_2_387 (.ZN (n_0_2_241), .A1 (n_0_2_240), .A2 (sps__n1), .B1 (n_0_2_234), .B2 (sps__n7));
OAI22_X1 i_0_2_386 (.ZN (n_0_2_240), .A1 (n_0_2_227), .A2 (n_0_2_154), .B1 (sps__n4), .B2 (n_0_2_239));
OAI221_X1 i_0_2_385 (.ZN (n_0_2_239), .A (n_0_2_208), .B1 (\multiplicand1[15] ), .B2 (spc__n22)
    , .C1 (spc__n19), .C2 (\multiplicand1[7] ));
OAI22_X1 i_0_2_384 (.ZN (n_0_274), .A1 (n_0_2_238), .A2 (sps__n10), .B1 (n_0_2_235), .B2 (n_0_2_148));
AOI22_X1 i_0_2_383 (.ZN (n_0_2_238), .A1 (n_0_2_237), .A2 (sps__n1), .B1 (n_0_2_231), .B2 (sps__n7));
OAI22_X1 i_0_2_382 (.ZN (n_0_2_237), .A1 (n_0_2_221), .A2 (n_0_2_154), .B1 (sps__n4), .B2 (n_0_2_236));
OAI221_X1 i_0_2_381 (.ZN (n_0_2_236), .A (n_0_2_208), .B1 (\multiplicand1[14] ), .B2 (spc__n22)
    , .C1 (spc__n19), .C2 (\multiplicand1[6] ));
OAI22_X1 i_0_2_380 (.ZN (n_0_273), .A1 (n_0_2_235), .A2 (sps__n10), .B1 (n_0_2_232), .B2 (n_0_2_148));
AOI22_X1 i_0_2_379 (.ZN (n_0_2_235), .A1 (n_0_2_228), .A2 (sps__n7), .B1 (n_0_2_234), .B2 (sps__n1));
OAI22_X1 i_0_2_378 (.ZN (n_0_2_234), .A1 (n_0_2_233), .A2 (sps__n4), .B1 (n_0_2_213), .B2 (n_0_2_154));
OAI221_X1 i_0_2_377 (.ZN (n_0_2_233), .A (n_0_2_208), .B1 (\multiplicand1[13] ), .B2 (spc__n22)
    , .C1 (spc__n19), .C2 (\multiplicand1[5] ));
OAI22_X1 i_0_2_376 (.ZN (n_0_272), .A1 (n_0_2_232), .A2 (sps__n10), .B1 (n_0_2_229), .B2 (n_0_2_148));
AOI22_X1 i_0_2_375 (.ZN (n_0_2_232), .A1 (n_0_2_222), .A2 (sps__n7), .B1 (n_0_2_231), .B2 (sps__n1));
OAI22_X1 i_0_2_374 (.ZN (n_0_2_231), .A1 (n_0_2_209), .A2 (n_0_2_154), .B1 (n_0_2_230), .B2 (sps__n4));
OAI221_X1 i_0_2_373 (.ZN (n_0_2_230), .A (n_0_2_208), .B1 (\multiplicand1[12] ), .B2 (spc__n22)
    , .C1 (spc__n19), .C2 (\multiplicand1[4] ));
OAI22_X1 i_0_2_372 (.ZN (n_0_271), .A1 (n_0_2_229), .A2 (sps__n10), .B1 (n_0_2_223), .B2 (n_0_2_148));
AOI22_X1 i_0_2_371 (.ZN (n_0_2_229), .A1 (n_0_2_228), .A2 (sps__n1), .B1 (sps__n7), .B2 (n_0_2_214));
OAI21_X1 i_0_2_370 (.ZN (n_0_2_228), .A (n_0_2_224), .B1 (n_0_2_227), .B2 (sps__n4));
INV_X1 i_0_2_369 (.ZN (n_0_2_227), .A (n_0_2_226));
OAI33_X1 i_0_2_368 (.ZN (n_0_2_226), .A1 (n_0_2_217), .A2 (n_0_2_225), .A3 (spc__n22)
    , .B1 (n_0_2_219), .B2 (spc__n16), .B3 (n_0_2_203));
INV_X1 i_0_2_367 (.ZN (n_0_2_225), .A (\multiplicand1[11] ));
NAND3_X1 i_0_2_366 (.ZN (n_0_2_224), .A1 (n_0_2_181), .A2 (\multiplicand1[7] ), .A3 (sps__n4));
OAI22_X1 i_0_2_365 (.ZN (n_0_270), .A1 (n_0_2_223), .A2 (sps__n10), .B1 (n_0_2_148), .B2 (n_0_2_215));
AOI22_X1 i_0_2_364 (.ZN (n_0_2_223), .A1 (n_0_2_222), .A2 (sps__n1), .B1 (sps__n7), .B2 (n_0_2_210));
OAI21_X1 i_0_2_363 (.ZN (n_0_2_222), .A (n_0_2_216), .B1 (n_0_2_221), .B2 (sps__n4));
INV_X1 i_0_2_362 (.ZN (n_0_2_221), .A (n_0_2_220));
OAI33_X1 i_0_2_361 (.ZN (n_0_2_220), .A1 (n_0_2_217), .A2 (n_0_2_218), .A3 (spc__n22)
    , .B1 (n_0_2_219), .B2 (spc__n16), .B3 (n_0_2_198));
NAND2_X1 i_0_2_360 (.ZN (n_0_2_219), .A1 (n_0_2_10), .A2 (spc__n22));
INV_X1 i_0_2_359 (.ZN (n_0_2_218), .A (\multiplicand1[10] ));
INV_X1 i_0_2_358 (.ZN (n_0_2_217), .A (n_0_2_208));
NAND3_X1 i_0_2_357 (.ZN (n_0_2_216), .A1 (n_0_2_181), .A2 (\multiplicand1[6] ), .A3 (sps__n4));
OAI22_X1 i_0_2_356 (.ZN (n_0_269), .A1 (n_0_2_215), .A2 (sps__n10), .B1 (n_0_2_211), .B2 (n_0_2_148));
AOI22_X1 i_0_2_355 (.ZN (n_0_2_215), .A1 (n_0_2_214), .A2 (sps__n1), .B1 (n_0_2_205), .B2 (sps__n7));
OAI21_X1 i_0_2_354 (.ZN (n_0_2_214), .A (n_0_2_212), .B1 (n_0_2_213), .B2 (sps__n4));
OAI221_X1 i_0_2_353 (.ZN (n_0_2_213), .A (n_0_2_208), .B1 (\multiplicand1[9] ), .B2 (spc__n22)
    , .C1 (spc__n19), .C2 (\multiplicand1[1] ));
NAND3_X1 i_0_2_352 (.ZN (n_0_2_212), .A1 (n_0_2_181), .A2 (\multiplicand1[5] ), .A3 (sps__n4));
OAI22_X1 i_0_2_351 (.ZN (n_0_268), .A1 (n_0_2_211), .A2 (sps__n10), .B1 (n_0_2_206), .B2 (n_0_2_148));
AOI22_X1 i_0_2_350 (.ZN (n_0_2_211), .A1 (n_0_2_210), .A2 (sps__n1), .B1 (n_0_2_200), .B2 (sps__n7));
OAI21_X1 i_0_2_349 (.ZN (n_0_2_210), .A (n_0_2_207), .B1 (n_0_2_209), .B2 (sps__n4));
OAI221_X1 i_0_2_348 (.ZN (n_0_2_209), .A (n_0_2_208), .B1 (\multiplicand1[8] ), .B2 (spc__n22)
    , .C1 (spc__n19), .C2 (\multiplicand1[0] ));
NOR2_X1 i_0_2_347 (.ZN (n_0_2_208), .A1 (spc__n16), .A2 (\counter[5] ));
NAND3_X1 i_0_2_346 (.ZN (n_0_2_207), .A1 (n_0_2_181), .A2 (\multiplicand1[4] ), .A3 (sps__n4));
OAI22_X1 i_0_2_345 (.ZN (n_0_267), .A1 (n_0_2_202), .A2 (n_0_2_148), .B1 (n_0_2_206), .B2 (sps__n10));
AOI22_X1 i_0_2_344 (.ZN (n_0_2_206), .A1 (n_0_2_205), .A2 (sps__n1), .B1 (n_0_2_196), .B2 (n_0_2_201));
AOI221_X1 i_0_2_343 (.ZN (n_0_2_205), .A (n_0_2_182), .B1 (n_0_2_203), .B2 (sps__n4)
    , .C1 (n_0_2_204), .C2 (n_0_2_154));
INV_X1 i_0_2_342 (.ZN (n_0_2_204), .A (\multiplicand1[7] ));
INV_X1 i_0_2_341 (.ZN (n_0_2_203), .A (\multiplicand1[3] ));
OAI22_X1 i_0_2_340 (.ZN (n_0_266), .A1 (n_0_2_202), .A2 (sps__n10), .B1 (n_0_2_194), .B2 (n_0_2_197));
AOI22_X1 i_0_2_339 (.ZN (n_0_2_202), .A1 (n_0_2_200), .A2 (sps__n1), .B1 (n_0_2_191), .B2 (n_0_2_201));
NOR2_X1 i_0_2_338 (.ZN (n_0_2_201), .A1 (n_0_2_182), .A2 (sps__n1));
AOI221_X1 i_0_2_337 (.ZN (n_0_2_200), .A (n_0_2_182), .B1 (n_0_2_198), .B2 (sps__n4)
    , .C1 (n_0_2_199), .C2 (n_0_2_154));
INV_X1 i_0_2_336 (.ZN (n_0_2_199), .A (\multiplicand1[6] ));
INV_X1 i_0_2_335 (.ZN (n_0_2_198), .A (\multiplicand1[2] ));
OAI33_X1 i_0_2_334 (.ZN (n_0_265), .A1 (n_0_2_197), .A2 (sps__n10), .A3 (n_0_2_182)
    , .B1 (n_0_2_193), .B2 (n_0_2_148), .B3 (n_0_2_182));
AOI22_X1 i_0_2_333 (.ZN (n_0_2_197), .A1 (n_0_2_196), .A2 (sps__n1), .B1 (n_0_2_192), .B2 (\multiplicand1[3] ));
OAI22_X1 i_0_2_332 (.ZN (n_0_2_196), .A1 (n_0_2_185), .A2 (n_0_2_154), .B1 (n_0_2_195), .B2 (sps__n4));
INV_X1 i_0_2_331 (.ZN (n_0_2_195), .A (\multiplicand1[5] ));
OAI33_X1 i_0_2_330 (.ZN (n_0_264), .A1 (n_0_2_193), .A2 (sps__n10), .A3 (n_0_2_182)
    , .B1 (n_0_2_194), .B2 (sps__n4), .B3 (n_0_2_189));
NAND2_X1 i_0_2_329 (.ZN (n_0_2_194), .A1 (n_0_2_181), .A2 (sps__n10));
AOI22_X1 i_0_2_328 (.ZN (n_0_2_193), .A1 (n_0_2_191), .A2 (sps__n1), .B1 (n_0_2_192), .B2 (\multiplicand1[2] ));
INV_X1 i_0_2_327 (.ZN (n_0_2_192), .A (n_0_2_155));
OAI22_X1 i_0_2_326 (.ZN (n_0_2_191), .A1 (n_0_2_183), .A2 (n_0_2_154), .B1 (n_0_2_190), .B2 (sps__n4));
INV_X1 i_0_2_325 (.ZN (n_0_2_190), .A (\multiplicand1[4] ));
AOI221_X1 i_0_2_324 (.ZN (n_0_263), .A (n_0_2_186), .B1 (n_0_2_188), .B2 (sps__n10)
    , .C1 (n_0_2_148), .C2 (n_0_2_189));
AOI22_X1 i_0_2_323 (.ZN (n_0_2_189), .A1 (sps__n1), .A2 (\multiplicand1[3] ), .B1 (\multiplicand1[1] ), .B2 (sps__n7));
AOI221_X1 i_0_2_322 (.ZN (n_0_262), .A (n_0_2_186), .B1 (sps__n10), .B2 (n_0_2_187)
    , .C1 (n_0_2_188), .C2 (n_0_2_148));
AOI22_X1 i_0_2_321 (.ZN (n_0_2_188), .A1 (sps__n1), .A2 (\multiplicand1[2] ), .B1 (\multiplicand1[0] ), .B2 (sps__n7));
NAND2_X1 i_0_2_320 (.ZN (n_0_2_187), .A1 (sps__n1), .A2 (\multiplicand1[1] ));
NAND2_X1 i_0_2_319 (.ZN (n_0_2_186), .A1 (n_0_2_181), .A2 (n_0_2_154));
AOI221_X1 i_0_2_318 (.ZN (n_0_261), .A (n_0_2_184), .B1 (n_0_2_183), .B2 (sps__n10)
    , .C1 (n_0_2_185), .C2 (n_0_2_148));
INV_X1 i_0_2_317 (.ZN (n_0_2_185), .A (\multiplicand1[1] ));
NAND2_X1 i_0_2_316 (.ZN (n_0_2_184), .A1 (n_0_2_181), .A2 (n_0_2_11));
NOR4_X1 i_0_2_315 (.ZN (n_0_260), .A1 (n_0_2_182), .A2 (n_0_2_12), .A3 (n_0_2_183), .A4 (sps__n10));
INV_X1 i_0_2_314 (.ZN (n_0_2_183), .A (\multiplicand1[0] ));
INV_X1 i_0_2_313 (.ZN (n_0_2_182), .A (n_0_2_181));
AND2_X1 i_0_2_312 (.ZN (n_0_2_181), .A1 (n_0_2_180), .A2 (n_0_2_13));
NOR2_X1 i_0_2_311 (.ZN (n_0_2_180), .A1 (\counter[5] ), .A2 (spc__n22));
OAI211_X1 i_0_2_310 (.ZN (n_0_389), .A (n_0_2_167), .B (n_0_2_16), .C1 (spc__n16), .C2 (n_0_2_179));
NAND2_X1 i_0_2_309 (.ZN (n_0_2_179), .A1 (n_0_2_172), .A2 (n_0_2_178));
OAI211_X1 i_0_2_308 (.ZN (n_0_2_178), .A (n_0_2_175), .B (spc__n19), .C1 (n_0_2_176), .C2 (n_0_2_177));
OAI22_X1 i_0_2_307 (.ZN (n_0_2_177), .A1 (n_0_2_12), .A2 (\multiplier1[0] ), .B1 (n_0_2_150), .B2 (\multiplier1[4] ));
OAI221_X1 i_0_2_306 (.ZN (n_0_2_176), .A (spw__n323), .B1 (n_0_2_153), .B2 (\multiplier1[6] )
    , .C1 (n_0_2_155), .C2 (\multiplier1[2] ));
OR3_X1 i_0_2_305 (.ZN (n_0_2_175), .A1 (n_0_2_173), .A2 (n_0_2_174), .A3 (spw__n323));
OAI22_X1 i_0_2_304 (.ZN (n_0_2_174), .A1 (n_0_2_155), .A2 (\multiplier1[3] ), .B1 (n_0_2_153), .B2 (\multiplier1[7] ));
OAI22_X1 i_0_2_303 (.ZN (n_0_2_173), .A1 (n_0_2_12), .A2 (\multiplier1[1] ), .B1 (n_0_2_150), .B2 (\multiplier1[5] ));
OAI221_X1 i_0_2_302 (.ZN (n_0_2_172), .A (spc__n22), .B1 (n_0_2_168), .B2 (n_0_2_169)
    , .C1 (n_0_2_170), .C2 (n_0_2_171));
OAI21_X1 i_0_2_301 (.ZN (n_0_2_171), .A (sps__n10), .B1 (n_0_2_155), .B2 (\multiplier1[11] ));
OAI222_X1 i_0_2_300 (.ZN (n_0_2_170), .A1 (n_0_2_12), .A2 (\multiplier1[9] ), .B1 (n_0_2_150)
    , .B2 (\multiplier1[13] ), .C1 (n_0_2_153), .C2 (\multiplier1[15] ));
OAI22_X1 i_0_2_299 (.ZN (n_0_2_169), .A1 (n_0_2_12), .A2 (\multiplier1[8] ), .B1 (n_0_2_155), .B2 (\multiplier1[10] ));
OAI221_X1 i_0_2_298 (.ZN (n_0_2_168), .A (spw__n323), .B1 (n_0_2_153), .B2 (\multiplier1[14] )
    , .C1 (n_0_2_150), .C2 (\multiplier1[12] ));
AOI21_X1 i_0_2_297 (.ZN (n_0_2_167), .A (n_0_2_160), .B1 (n_0_2_161), .B2 (n_0_2_166));
OAI22_X1 i_0_2_296 (.ZN (n_0_2_166), .A1 (n_0_2_162), .A2 (n_0_2_163), .B1 (n_0_2_164), .B2 (n_0_2_165));
OAI22_X1 i_0_2_295 (.ZN (n_0_2_165), .A1 (n_0_2_12), .A2 (\multiplier1[16] ), .B1 (n_0_2_153), .B2 (\multiplier1[22] ));
OAI221_X1 i_0_2_294 (.ZN (n_0_2_164), .A (spw__n323), .B1 (n_0_2_155), .B2 (\multiplier1[18] )
    , .C1 (\multiplier1[20] ), .C2 (n_0_2_150));
OAI21_X1 i_0_2_293 (.ZN (n_0_2_163), .A (sps__n10), .B1 (n_0_2_155), .B2 (\multiplier1[19] ));
OAI222_X1 i_0_2_292 (.ZN (n_0_2_162), .A1 (n_0_2_12), .A2 (\multiplier1[17] ), .B1 (n_0_2_150)
    , .B2 (\multiplier1[21] ), .C1 (n_0_2_153), .C2 (\multiplier1[23] ));
NOR2_X1 i_0_2_291 (.ZN (n_0_2_161), .A1 (n_0_2_13), .A2 (spc__n22));
AOI211_X1 i_0_2_290 (.ZN (n_0_2_160), .A (n_0_2_13), .B (spc__n19), .C1 (n_0_2_156), .C2 (n_0_2_159));
OAI221_X1 i_0_2_289 (.ZN (n_0_2_159), .A (n_0_2_158), .B1 (\multiplier1[29] ), .B2 (n_0_2_150)
    , .C1 (\multiplier1[25] ), .C2 (n_0_2_12));
INV_X1 i_0_2_288 (.ZN (n_0_2_158), .A (n_0_2_157));
OAI221_X1 i_0_2_287 (.ZN (n_0_2_157), .A (sps__n10), .B1 (n_0_2_153), .B2 (\multiplier1[31] )
    , .C1 (n_0_2_155), .C2 (\multiplier1[27] ));
OAI221_X1 i_0_2_286 (.ZN (n_0_2_156), .A (n_0_2_152), .B1 (\multiplier1[30] ), .B2 (n_0_2_153)
    , .C1 (\multiplier1[26] ), .C2 (n_0_2_155));
NAND2_X4 i_0_2_285 (.ZN (n_0_2_155), .A1 (n_0_2_154), .A2 (sps__n7));
INV_X32 i_0_2_284 (.ZN (n_0_2_154), .A (sps__n4));
NAND2_X1 i_0_2_283 (.ZN (n_0_2_153), .A1 (sps__n4), .A2 (sps__n7));
INV_X1 i_0_2_282 (.ZN (n_0_2_152), .A (n_0_2_151));
OAI221_X1 i_0_2_281 (.ZN (n_0_2_151), .A (spw__n323), .B1 (n_0_2_150), .B2 (\multiplier1[28] )
    , .C1 (n_0_2_12), .C2 (\multiplier1[24] ));
NAND2_X2 i_0_2_280 (.ZN (n_0_2_150), .A1 (sps__n1), .A2 (sps__n4));
INV_X4 i_0_2_279 (.ZN (n_0_2_149), .A (sps__n7));
INV_X4 i_0_2_278 (.ZN (n_0_2_148), .A (sps__n10));
INV_X1 i_0_2_277 (.ZN (n_0_2_147), .A (spc__n22));
OAI22_X1 i_0_2_276 (.ZN (n_0_388), .A1 (n_0_2_20), .A2 (n_0_2_145), .B1 (n_0_2_21), .B2 (n_0_2_146));
INV_X1 i_0_2_275 (.ZN (n_0_2_146), .A (n_0_190));
INV_X1 i_0_2_274 (.ZN (n_0_452), .A (n_0_2_145));
AOI22_X1 i_0_2_273 (.ZN (n_0_2_145), .A1 (n_0_2_18), .A2 (\accumulator[63] ), .B1 (n_0_64), .B2 (sps__n13));
OAI22_X1 i_0_2_272 (.ZN (n_0_387), .A1 (n_0_2_20), .A2 (n_0_2_143), .B1 (n_0_2_21), .B2 (n_0_2_144));
INV_X1 i_0_2_271 (.ZN (n_0_2_144), .A (n_0_189));
INV_X1 i_0_2_270 (.ZN (n_0_451), .A (n_0_2_143));
AOI22_X1 i_0_2_269 (.ZN (n_0_2_143), .A1 (n_0_2_18), .A2 (\accumulator[62] ), .B1 (n_0_63), .B2 (sps__n13));
OAI22_X1 i_0_2_268 (.ZN (n_0_386), .A1 (n_0_2_20), .A2 (n_0_2_141), .B1 (n_0_2_21), .B2 (n_0_2_142));
INV_X1 i_0_2_267 (.ZN (n_0_2_142), .A (n_0_188));
INV_X1 i_0_2_266 (.ZN (n_0_450), .A (n_0_2_141));
AOI22_X2 i_0_2_265 (.ZN (n_0_2_141), .A1 (n_0_2_18), .A2 (\accumulator[61] ), .B1 (n_0_62), .B2 (sps__n13));
OAI22_X1 i_0_2_264 (.ZN (n_0_385), .A1 (n_0_2_20), .A2 (n_0_2_139), .B1 (n_0_2_21), .B2 (n_0_2_140));
INV_X1 i_0_2_263 (.ZN (n_0_2_140), .A (n_0_187));
INV_X1 i_0_2_262 (.ZN (n_0_449), .A (n_0_2_139));
AOI22_X1 i_0_2_261 (.ZN (n_0_2_139), .A1 (n_0_2_18), .A2 (\accumulator[60] ), .B1 (n_0_61), .B2 (sps__n13));
OAI22_X1 i_0_2_260 (.ZN (n_0_384), .A1 (n_0_2_20), .A2 (n_0_2_137), .B1 (n_0_2_21), .B2 (n_0_2_138));
INV_X1 i_0_2_259 (.ZN (n_0_2_138), .A (n_0_186));
INV_X1 i_0_2_258 (.ZN (n_0_448), .A (n_0_2_137));
AOI22_X1 i_0_2_257 (.ZN (n_0_2_137), .A1 (n_0_2_18), .A2 (\accumulator[59] ), .B1 (n_0_60), .B2 (sps__n13));
OAI22_X1 i_0_2_256 (.ZN (n_0_383), .A1 (n_0_2_20), .A2 (n_0_2_135), .B1 (n_0_2_21), .B2 (n_0_2_136));
INV_X1 i_0_2_255 (.ZN (n_0_2_136), .A (n_0_185));
INV_X1 i_0_2_254 (.ZN (n_0_447), .A (n_0_2_135));
AOI22_X1 i_0_2_253 (.ZN (n_0_2_135), .A1 (n_0_2_18), .A2 (\accumulator[58] ), .B1 (n_0_59), .B2 (sps__n13));
OAI22_X1 i_0_2_252 (.ZN (n_0_382), .A1 (n_0_2_20), .A2 (n_0_2_133), .B1 (n_0_2_21), .B2 (n_0_2_134));
INV_X1 i_0_2_251 (.ZN (n_0_2_134), .A (n_0_184));
INV_X1 i_0_2_250 (.ZN (n_0_446), .A (n_0_2_133));
AOI22_X1 i_0_2_249 (.ZN (n_0_2_133), .A1 (n_0_2_18), .A2 (\accumulator[57] ), .B1 (n_0_58), .B2 (sps__n13));
OAI22_X1 i_0_2_248 (.ZN (n_0_381), .A1 (n_0_2_20), .A2 (n_0_2_131), .B1 (n_0_2_21), .B2 (n_0_2_132));
INV_X1 i_0_2_247 (.ZN (n_0_2_132), .A (n_0_183));
INV_X1 i_0_2_246 (.ZN (n_0_445), .A (n_0_2_131));
AOI22_X1 i_0_2_245 (.ZN (n_0_2_131), .A1 (n_0_2_18), .A2 (\accumulator[56] ), .B1 (n_0_57), .B2 (sps__n13));
OAI22_X1 i_0_2_244 (.ZN (n_0_380), .A1 (n_0_2_20), .A2 (n_0_2_129), .B1 (n_0_2_21), .B2 (n_0_2_130));
INV_X1 i_0_2_243 (.ZN (n_0_2_130), .A (n_0_182));
INV_X1 i_0_2_242 (.ZN (n_0_444), .A (n_0_2_129));
AOI22_X1 i_0_2_241 (.ZN (n_0_2_129), .A1 (n_0_2_18), .A2 (\accumulator[55] ), .B1 (n_0_56), .B2 (sps__n13));
OAI22_X1 i_0_2_240 (.ZN (n_0_379), .A1 (n_0_2_20), .A2 (n_0_2_127), .B1 (n_0_2_21), .B2 (n_0_2_128));
INV_X1 i_0_2_239 (.ZN (n_0_2_128), .A (n_0_181));
INV_X1 i_0_2_238 (.ZN (n_0_443), .A (n_0_2_127));
AOI22_X1 i_0_2_237 (.ZN (n_0_2_127), .A1 (n_0_2_18), .A2 (\accumulator[54] ), .B1 (n_0_55), .B2 (sps__n13));
OAI22_X1 i_0_2_236 (.ZN (n_0_378), .A1 (n_0_2_20), .A2 (n_0_2_125), .B1 (n_0_2_21), .B2 (n_0_2_126));
INV_X1 i_0_2_235 (.ZN (n_0_2_126), .A (n_0_180));
INV_X1 i_0_2_234 (.ZN (n_0_442), .A (n_0_2_125));
AOI22_X1 i_0_2_233 (.ZN (n_0_2_125), .A1 (n_0_2_18), .A2 (\accumulator[53] ), .B1 (n_0_54), .B2 (sps__n13));
OAI22_X1 i_0_2_232 (.ZN (n_0_377), .A1 (n_0_2_20), .A2 (n_0_2_123), .B1 (n_0_2_21), .B2 (n_0_2_124));
INV_X1 i_0_2_231 (.ZN (n_0_2_124), .A (n_0_179));
INV_X1 i_0_2_230 (.ZN (n_0_441), .A (n_0_2_123));
AOI22_X1 i_0_2_229 (.ZN (n_0_2_123), .A1 (n_0_2_18), .A2 (\accumulator[52] ), .B1 (n_0_53), .B2 (sps__n13));
OAI22_X1 i_0_2_228 (.ZN (n_0_376), .A1 (n_0_2_20), .A2 (n_0_2_121), .B1 (n_0_2_21), .B2 (n_0_2_122));
INV_X1 i_0_2_227 (.ZN (n_0_2_122), .A (n_0_178));
INV_X1 i_0_2_226 (.ZN (n_0_440), .A (n_0_2_121));
AOI22_X1 i_0_2_225 (.ZN (n_0_2_121), .A1 (n_0_2_18), .A2 (\accumulator[51] ), .B1 (n_0_52), .B2 (sps__n13));
OAI22_X1 i_0_2_224 (.ZN (n_0_375), .A1 (n_0_2_20), .A2 (n_0_2_119), .B1 (n_0_2_21), .B2 (n_0_2_120));
INV_X1 i_0_2_223 (.ZN (n_0_2_120), .A (n_0_177));
INV_X1 i_0_2_222 (.ZN (n_0_439), .A (n_0_2_119));
AOI22_X1 i_0_2_221 (.ZN (n_0_2_119), .A1 (n_0_2_18), .A2 (\accumulator[50] ), .B1 (n_0_51), .B2 (sps__n13));
OAI22_X1 i_0_2_220 (.ZN (n_0_374), .A1 (n_0_2_20), .A2 (n_0_2_117), .B1 (n_0_2_21), .B2 (n_0_2_118));
INV_X1 i_0_2_219 (.ZN (n_0_2_118), .A (n_0_176));
INV_X1 i_0_2_218 (.ZN (n_0_438), .A (n_0_2_117));
AOI22_X1 i_0_2_217 (.ZN (n_0_2_117), .A1 (n_0_2_18), .A2 (\accumulator[49] ), .B1 (n_0_50), .B2 (sps__n13));
OAI22_X1 i_0_2_216 (.ZN (n_0_373), .A1 (n_0_2_20), .A2 (n_0_2_115), .B1 (n_0_2_21), .B2 (n_0_2_116));
INV_X1 i_0_2_215 (.ZN (n_0_2_116), .A (n_0_175));
INV_X1 i_0_2_214 (.ZN (n_0_437), .A (n_0_2_115));
AOI22_X1 i_0_2_213 (.ZN (n_0_2_115), .A1 (n_0_2_18), .A2 (\accumulator[48] ), .B1 (n_0_49), .B2 (sps__n13));
OAI22_X1 i_0_2_212 (.ZN (n_0_372), .A1 (n_0_2_20), .A2 (n_0_2_113), .B1 (n_0_2_21), .B2 (n_0_2_114));
INV_X1 i_0_2_211 (.ZN (n_0_2_114), .A (n_0_174));
INV_X1 i_0_2_210 (.ZN (n_0_436), .A (n_0_2_113));
AOI22_X1 i_0_2_209 (.ZN (n_0_2_113), .A1 (n_0_2_18), .A2 (\accumulator[47] ), .B1 (n_0_48), .B2 (sps__n13));
OAI22_X1 i_0_2_208 (.ZN (n_0_371), .A1 (n_0_2_20), .A2 (n_0_2_111), .B1 (n_0_2_21), .B2 (n_0_2_112));
INV_X1 i_0_2_207 (.ZN (n_0_2_112), .A (n_0_173));
INV_X1 i_0_2_206 (.ZN (n_0_435), .A (n_0_2_111));
AOI22_X1 i_0_2_205 (.ZN (n_0_2_111), .A1 (n_0_2_18), .A2 (\accumulator[46] ), .B1 (n_0_47), .B2 (sps__n13));
OAI22_X1 i_0_2_204 (.ZN (n_0_370), .A1 (n_0_2_20), .A2 (n_0_2_109), .B1 (n_0_2_21), .B2 (n_0_2_110));
INV_X1 i_0_2_203 (.ZN (n_0_2_110), .A (n_0_172));
INV_X1 i_0_2_202 (.ZN (n_0_434), .A (n_0_2_109));
AOI22_X1 i_0_2_201 (.ZN (n_0_2_109), .A1 (n_0_2_18), .A2 (\accumulator[45] ), .B1 (n_0_46), .B2 (sps__n13));
OAI22_X1 i_0_2_200 (.ZN (n_0_369), .A1 (n_0_2_20), .A2 (n_0_2_107), .B1 (n_0_2_21), .B2 (n_0_2_108));
INV_X1 i_0_2_199 (.ZN (n_0_2_108), .A (n_0_171));
INV_X1 i_0_2_198 (.ZN (n_0_433), .A (n_0_2_107));
AOI22_X1 i_0_2_197 (.ZN (n_0_2_107), .A1 (n_0_2_18), .A2 (\accumulator[44] ), .B1 (n_0_45), .B2 (sps__n13));
OAI22_X1 i_0_2_196 (.ZN (n_0_368), .A1 (n_0_2_20), .A2 (n_0_2_105), .B1 (n_0_2_21), .B2 (n_0_2_106));
INV_X1 i_0_2_195 (.ZN (n_0_2_106), .A (n_0_170));
INV_X1 i_0_2_194 (.ZN (n_0_432), .A (n_0_2_105));
AOI22_X1 i_0_2_193 (.ZN (n_0_2_105), .A1 (n_0_2_18), .A2 (\accumulator[43] ), .B1 (n_0_44), .B2 (sps__n13));
OAI22_X1 i_0_2_192 (.ZN (n_0_367), .A1 (n_0_2_20), .A2 (n_0_2_103), .B1 (n_0_2_21), .B2 (n_0_2_104));
INV_X1 i_0_2_191 (.ZN (n_0_2_104), .A (n_0_169));
INV_X1 i_0_2_190 (.ZN (n_0_431), .A (n_0_2_103));
AOI22_X1 i_0_2_189 (.ZN (n_0_2_103), .A1 (n_0_2_18), .A2 (\accumulator[42] ), .B1 (n_0_43), .B2 (sps__n13));
OAI22_X1 i_0_2_188 (.ZN (n_0_366), .A1 (n_0_2_20), .A2 (n_0_2_101), .B1 (n_0_2_21), .B2 (n_0_2_102));
INV_X1 i_0_2_187 (.ZN (n_0_2_102), .A (n_0_168));
INV_X1 i_0_2_186 (.ZN (n_0_430), .A (n_0_2_101));
AOI22_X1 i_0_2_185 (.ZN (n_0_2_101), .A1 (n_0_2_18), .A2 (\accumulator[41] ), .B1 (n_0_42), .B2 (sps__n13));
OAI22_X1 i_0_2_184 (.ZN (n_0_365), .A1 (n_0_2_20), .A2 (n_0_2_99), .B1 (n_0_2_21), .B2 (n_0_2_100));
INV_X1 i_0_2_183 (.ZN (n_0_2_100), .A (n_0_167));
INV_X1 i_0_2_182 (.ZN (n_0_429), .A (n_0_2_99));
AOI22_X1 i_0_2_181 (.ZN (n_0_2_99), .A1 (n_0_2_18), .A2 (\accumulator[40] ), .B1 (n_0_41), .B2 (sps__n13));
OAI22_X1 i_0_2_180 (.ZN (n_0_364), .A1 (n_0_2_20), .A2 (n_0_2_97), .B1 (n_0_2_21), .B2 (n_0_2_98));
INV_X1 i_0_2_179 (.ZN (n_0_2_98), .A (n_0_166));
INV_X1 i_0_2_178 (.ZN (n_0_428), .A (n_0_2_97));
AOI22_X1 i_0_2_177 (.ZN (n_0_2_97), .A1 (n_0_2_18), .A2 (\accumulator[39] ), .B1 (n_0_40), .B2 (sps__n13));
OAI22_X1 i_0_2_176 (.ZN (n_0_363), .A1 (n_0_2_20), .A2 (n_0_2_95), .B1 (n_0_2_21), .B2 (n_0_2_96));
INV_X1 i_0_2_175 (.ZN (n_0_2_96), .A (n_0_165));
INV_X1 i_0_2_174 (.ZN (n_0_427), .A (n_0_2_95));
AOI22_X1 i_0_2_173 (.ZN (n_0_2_95), .A1 (n_0_2_18), .A2 (\accumulator[38] ), .B1 (n_0_39), .B2 (sps__n13));
OAI22_X1 i_0_2_172 (.ZN (n_0_362), .A1 (n_0_2_20), .A2 (n_0_2_93), .B1 (n_0_2_21), .B2 (n_0_2_94));
INV_X1 i_0_2_171 (.ZN (n_0_2_94), .A (n_0_164));
INV_X1 i_0_2_170 (.ZN (n_0_426), .A (n_0_2_93));
AOI22_X1 i_0_2_169 (.ZN (n_0_2_93), .A1 (n_0_2_18), .A2 (\accumulator[37] ), .B1 (n_0_38), .B2 (sps__n13));
OAI22_X1 i_0_2_168 (.ZN (n_0_361), .A1 (n_0_2_20), .A2 (n_0_2_91), .B1 (n_0_2_21), .B2 (n_0_2_92));
INV_X1 i_0_2_167 (.ZN (n_0_2_92), .A (n_0_163));
INV_X1 i_0_2_166 (.ZN (n_0_425), .A (n_0_2_91));
AOI22_X1 i_0_2_165 (.ZN (n_0_2_91), .A1 (n_0_2_18), .A2 (\accumulator[36] ), .B1 (n_0_37), .B2 (sps__n13));
OAI22_X1 i_0_2_164 (.ZN (n_0_360), .A1 (n_0_2_20), .A2 (n_0_2_89), .B1 (n_0_2_21), .B2 (n_0_2_90));
INV_X1 i_0_2_163 (.ZN (n_0_2_90), .A (n_0_162));
INV_X1 i_0_2_162 (.ZN (n_0_424), .A (n_0_2_89));
AOI22_X1 i_0_2_161 (.ZN (n_0_2_89), .A1 (n_0_2_18), .A2 (\accumulator[35] ), .B1 (n_0_36), .B2 (sps__n13));
OAI22_X1 i_0_2_160 (.ZN (n_0_359), .A1 (n_0_2_20), .A2 (n_0_2_87), .B1 (n_0_2_21), .B2 (n_0_2_88));
INV_X1 i_0_2_159 (.ZN (n_0_2_88), .A (n_0_161));
INV_X1 i_0_2_158 (.ZN (n_0_423), .A (n_0_2_87));
AOI22_X1 i_0_2_157 (.ZN (n_0_2_87), .A1 (n_0_2_18), .A2 (\accumulator[34] ), .B1 (n_0_35), .B2 (sps__n13));
OAI22_X1 i_0_2_156 (.ZN (n_0_358), .A1 (n_0_2_20), .A2 (n_0_2_85), .B1 (n_0_2_21), .B2 (n_0_2_86));
INV_X1 i_0_2_155 (.ZN (n_0_2_86), .A (n_0_160));
INV_X1 i_0_2_154 (.ZN (n_0_422), .A (n_0_2_85));
AOI22_X1 i_0_2_153 (.ZN (n_0_2_85), .A1 (n_0_2_18), .A2 (\accumulator[33] ), .B1 (n_0_34), .B2 (sps__n13));
OAI22_X1 i_0_2_152 (.ZN (n_0_357), .A1 (n_0_2_20), .A2 (n_0_2_83), .B1 (n_0_2_21), .B2 (n_0_2_84));
INV_X1 i_0_2_151 (.ZN (n_0_2_84), .A (n_0_159));
INV_X1 i_0_2_150 (.ZN (n_0_421), .A (n_0_2_83));
AOI22_X1 i_0_2_149 (.ZN (n_0_2_83), .A1 (n_0_2_18), .A2 (\accumulator[32] ), .B1 (n_0_33), .B2 (sps__n13));
OAI22_X1 i_0_2_148 (.ZN (n_0_356), .A1 (n_0_2_20), .A2 (n_0_2_81), .B1 (n_0_2_21), .B2 (n_0_2_82));
INV_X1 i_0_2_147 (.ZN (n_0_2_82), .A (n_0_158));
INV_X1 i_0_2_146 (.ZN (n_0_420), .A (n_0_2_81));
AOI22_X1 i_0_2_145 (.ZN (n_0_2_81), .A1 (n_0_2_18), .A2 (\accumulator[31] ), .B1 (n_0_32), .B2 (sps__n13));
OAI22_X1 i_0_2_144 (.ZN (n_0_355), .A1 (n_0_2_20), .A2 (n_0_2_79), .B1 (n_0_2_21), .B2 (n_0_2_80));
INV_X1 i_0_2_143 (.ZN (n_0_2_80), .A (n_0_157));
INV_X1 i_0_2_142 (.ZN (n_0_419), .A (n_0_2_79));
AOI22_X1 i_0_2_141 (.ZN (n_0_2_79), .A1 (n_0_2_18), .A2 (\accumulator[30] ), .B1 (n_0_31), .B2 (sps__n13));
OAI22_X1 i_0_2_140 (.ZN (n_0_354), .A1 (n_0_2_20), .A2 (n_0_2_77), .B1 (n_0_2_21), .B2 (n_0_2_78));
INV_X1 i_0_2_139 (.ZN (n_0_2_78), .A (n_0_156));
INV_X1 i_0_2_138 (.ZN (n_0_418), .A (n_0_2_77));
AOI22_X1 i_0_2_137 (.ZN (n_0_2_77), .A1 (n_0_2_18), .A2 (\accumulator[29] ), .B1 (n_0_30), .B2 (sps__n13));
OAI22_X1 i_0_2_136 (.ZN (n_0_353), .A1 (n_0_2_20), .A2 (n_0_2_75), .B1 (n_0_2_21), .B2 (n_0_2_76));
INV_X1 i_0_2_135 (.ZN (n_0_2_76), .A (n_0_155));
INV_X1 i_0_2_134 (.ZN (n_0_417), .A (n_0_2_75));
AOI22_X1 i_0_2_133 (.ZN (n_0_2_75), .A1 (n_0_2_18), .A2 (\accumulator[28] ), .B1 (n_0_29), .B2 (sps__n13));
OAI22_X1 i_0_2_132 (.ZN (n_0_352), .A1 (n_0_2_20), .A2 (n_0_2_73), .B1 (n_0_2_21), .B2 (n_0_2_74));
INV_X1 i_0_2_131 (.ZN (n_0_2_74), .A (n_0_154));
INV_X1 i_0_2_130 (.ZN (n_0_416), .A (n_0_2_73));
AOI22_X1 i_0_2_129 (.ZN (n_0_2_73), .A1 (n_0_2_18), .A2 (\accumulator[27] ), .B1 (n_0_28), .B2 (sps__n13));
OAI22_X1 i_0_2_128 (.ZN (n_0_351), .A1 (n_0_2_20), .A2 (n_0_2_71), .B1 (n_0_2_21), .B2 (n_0_2_72));
INV_X1 i_0_2_127 (.ZN (n_0_2_72), .A (n_0_153));
INV_X1 i_0_2_126 (.ZN (n_0_415), .A (n_0_2_71));
AOI22_X1 i_0_2_125 (.ZN (n_0_2_71), .A1 (n_0_2_18), .A2 (\accumulator[26] ), .B1 (n_0_27), .B2 (sps__n13));
OAI22_X1 i_0_2_124 (.ZN (n_0_350), .A1 (n_0_2_20), .A2 (n_0_2_69), .B1 (n_0_2_21), .B2 (n_0_2_70));
INV_X1 i_0_2_123 (.ZN (n_0_2_70), .A (n_0_152));
INV_X1 i_0_2_122 (.ZN (n_0_414), .A (n_0_2_69));
AOI22_X1 i_0_2_121 (.ZN (n_0_2_69), .A1 (n_0_2_18), .A2 (\accumulator[25] ), .B1 (n_0_26), .B2 (sps__n13));
OAI22_X1 i_0_2_120 (.ZN (n_0_349), .A1 (n_0_2_20), .A2 (n_0_2_67), .B1 (n_0_2_21), .B2 (n_0_2_68));
INV_X1 i_0_2_119 (.ZN (n_0_2_68), .A (n_0_151));
INV_X1 i_0_2_118 (.ZN (n_0_413), .A (n_0_2_67));
AOI22_X1 i_0_2_117 (.ZN (n_0_2_67), .A1 (n_0_2_18), .A2 (\accumulator[24] ), .B1 (n_0_25), .B2 (sps__n13));
OAI22_X1 i_0_2_116 (.ZN (n_0_348), .A1 (n_0_2_20), .A2 (n_0_2_65), .B1 (n_0_2_21), .B2 (n_0_2_66));
INV_X1 i_0_2_115 (.ZN (n_0_2_66), .A (n_0_150));
INV_X1 i_0_2_114 (.ZN (n_0_412), .A (n_0_2_65));
AOI22_X1 i_0_2_113 (.ZN (n_0_2_65), .A1 (n_0_2_18), .A2 (\accumulator[23] ), .B1 (n_0_24), .B2 (sps__n13));
OAI22_X1 i_0_2_112 (.ZN (n_0_347), .A1 (n_0_2_20), .A2 (n_0_2_63), .B1 (n_0_2_21), .B2 (n_0_2_64));
INV_X1 i_0_2_111 (.ZN (n_0_2_64), .A (n_0_149));
INV_X1 i_0_2_110 (.ZN (n_0_411), .A (n_0_2_63));
AOI22_X1 i_0_2_109 (.ZN (n_0_2_63), .A1 (n_0_2_18), .A2 (\accumulator[22] ), .B1 (n_0_23), .B2 (sps__n13));
OAI22_X1 i_0_2_108 (.ZN (n_0_346), .A1 (n_0_2_20), .A2 (n_0_2_61), .B1 (n_0_2_21), .B2 (n_0_2_62));
INV_X1 i_0_2_107 (.ZN (n_0_2_62), .A (n_0_148));
INV_X1 i_0_2_106 (.ZN (n_0_410), .A (n_0_2_61));
AOI22_X1 i_0_2_105 (.ZN (n_0_2_61), .A1 (n_0_2_18), .A2 (\accumulator[21] ), .B1 (n_0_22), .B2 (sps__n13));
OAI22_X1 i_0_2_104 (.ZN (n_0_345), .A1 (n_0_2_20), .A2 (n_0_2_59), .B1 (n_0_2_21), .B2 (n_0_2_60));
INV_X1 i_0_2_103 (.ZN (n_0_2_60), .A (n_0_147));
INV_X1 i_0_2_102 (.ZN (n_0_409), .A (n_0_2_59));
AOI22_X1 i_0_2_101 (.ZN (n_0_2_59), .A1 (n_0_2_18), .A2 (\accumulator[20] ), .B1 (n_0_21), .B2 (sps__n13));
OAI22_X1 i_0_2_100 (.ZN (n_0_344), .A1 (n_0_2_20), .A2 (n_0_2_57), .B1 (n_0_2_21), .B2 (n_0_2_58));
INV_X1 i_0_2_99 (.ZN (n_0_2_58), .A (n_0_146));
INV_X1 i_0_2_98 (.ZN (n_0_408), .A (n_0_2_57));
AOI22_X1 i_0_2_97 (.ZN (n_0_2_57), .A1 (n_0_2_18), .A2 (\accumulator[19] ), .B1 (n_0_20), .B2 (sps__n13));
OAI22_X1 i_0_2_96 (.ZN (n_0_343), .A1 (n_0_2_20), .A2 (n_0_2_55), .B1 (n_0_2_21), .B2 (n_0_2_56));
INV_X1 i_0_2_95 (.ZN (n_0_2_56), .A (n_0_145));
INV_X1 i_0_2_94 (.ZN (n_0_407), .A (n_0_2_55));
AOI22_X1 i_0_2_93 (.ZN (n_0_2_55), .A1 (n_0_2_18), .A2 (\accumulator[18] ), .B1 (n_0_19), .B2 (sps__n13));
OAI22_X1 i_0_2_92 (.ZN (n_0_342), .A1 (n_0_2_20), .A2 (n_0_2_53), .B1 (n_0_2_21), .B2 (n_0_2_54));
INV_X1 i_0_2_91 (.ZN (n_0_2_54), .A (n_0_144));
INV_X1 i_0_2_90 (.ZN (n_0_406), .A (n_0_2_53));
AOI22_X1 i_0_2_89 (.ZN (n_0_2_53), .A1 (n_0_2_18), .A2 (\accumulator[17] ), .B1 (n_0_18), .B2 (sps__n13));
OAI22_X1 i_0_2_88 (.ZN (n_0_341), .A1 (n_0_2_20), .A2 (n_0_2_51), .B1 (n_0_2_21), .B2 (n_0_2_52));
INV_X1 i_0_2_87 (.ZN (n_0_2_52), .A (n_0_143));
INV_X1 i_0_2_86 (.ZN (n_0_405), .A (n_0_2_51));
AOI22_X1 i_0_2_85 (.ZN (n_0_2_51), .A1 (n_0_2_18), .A2 (\accumulator[16] ), .B1 (n_0_17), .B2 (sps__n13));
OAI22_X1 i_0_2_84 (.ZN (n_0_340), .A1 (n_0_2_20), .A2 (n_0_2_49), .B1 (n_0_2_21), .B2 (n_0_2_50));
INV_X1 i_0_2_83 (.ZN (n_0_2_50), .A (n_0_142));
INV_X1 i_0_2_82 (.ZN (n_0_404), .A (n_0_2_49));
AOI22_X1 i_0_2_81 (.ZN (n_0_2_49), .A1 (n_0_2_18), .A2 (\accumulator[15] ), .B1 (n_0_16), .B2 (sps__n13));
OAI22_X1 i_0_2_80 (.ZN (n_0_339), .A1 (n_0_2_20), .A2 (n_0_2_47), .B1 (n_0_2_21), .B2 (n_0_2_48));
INV_X1 i_0_2_79 (.ZN (n_0_2_48), .A (n_0_141));
INV_X1 i_0_2_78 (.ZN (n_0_403), .A (n_0_2_47));
AOI22_X1 i_0_2_77 (.ZN (n_0_2_47), .A1 (n_0_2_18), .A2 (\accumulator[14] ), .B1 (n_0_15), .B2 (sps__n13));
OAI22_X1 i_0_2_76 (.ZN (n_0_338), .A1 (n_0_2_20), .A2 (n_0_2_45), .B1 (n_0_2_21), .B2 (n_0_2_46));
INV_X1 i_0_2_75 (.ZN (n_0_2_46), .A (n_0_140));
INV_X1 i_0_2_74 (.ZN (n_0_402), .A (n_0_2_45));
AOI22_X1 i_0_2_73 (.ZN (n_0_2_45), .A1 (n_0_2_18), .A2 (\accumulator[13] ), .B1 (n_0_14), .B2 (sps__n13));
OAI22_X1 i_0_2_72 (.ZN (n_0_337), .A1 (n_0_2_20), .A2 (n_0_2_43), .B1 (n_0_2_21), .B2 (n_0_2_44));
INV_X1 i_0_2_71 (.ZN (n_0_2_44), .A (n_0_139));
INV_X1 i_0_2_70 (.ZN (n_0_401), .A (n_0_2_43));
AOI22_X1 i_0_2_69 (.ZN (n_0_2_43), .A1 (n_0_2_18), .A2 (\accumulator[12] ), .B1 (n_0_13), .B2 (sps__n13));
OAI22_X1 i_0_2_68 (.ZN (n_0_336), .A1 (n_0_2_20), .A2 (n_0_2_41), .B1 (n_0_2_21), .B2 (n_0_2_42));
INV_X1 i_0_2_67 (.ZN (n_0_2_42), .A (n_0_138));
INV_X1 i_0_2_66 (.ZN (n_0_400), .A (n_0_2_41));
AOI22_X1 i_0_2_65 (.ZN (n_0_2_41), .A1 (n_0_2_18), .A2 (\accumulator[11] ), .B1 (n_0_12), .B2 (sps__n13));
OAI22_X1 i_0_2_64 (.ZN (n_0_335), .A1 (n_0_2_20), .A2 (n_0_2_39), .B1 (n_0_2_21), .B2 (n_0_2_40));
INV_X1 i_0_2_63 (.ZN (n_0_2_40), .A (n_0_137));
INV_X1 i_0_2_62 (.ZN (n_0_399), .A (n_0_2_39));
AOI22_X1 i_0_2_61 (.ZN (n_0_2_39), .A1 (n_0_2_18), .A2 (\accumulator[10] ), .B1 (n_0_11), .B2 (sps__n13));
OAI22_X1 i_0_2_60 (.ZN (n_0_334), .A1 (n_0_2_20), .A2 (n_0_2_37), .B1 (n_0_2_21), .B2 (n_0_2_38));
INV_X1 i_0_2_59 (.ZN (n_0_2_38), .A (n_0_136));
INV_X1 i_0_2_58 (.ZN (n_0_398), .A (n_0_2_37));
AOI22_X1 i_0_2_57 (.ZN (n_0_2_37), .A1 (n_0_2_18), .A2 (\accumulator[9] ), .B1 (n_0_10), .B2 (sps__n13));
OAI22_X1 i_0_2_56 (.ZN (n_0_333), .A1 (n_0_2_20), .A2 (n_0_2_35), .B1 (n_0_2_21), .B2 (n_0_2_36));
INV_X1 i_0_2_55 (.ZN (n_0_2_36), .A (n_0_135));
INV_X1 i_0_2_54 (.ZN (n_0_397), .A (n_0_2_35));
AOI22_X1 i_0_2_53 (.ZN (n_0_2_35), .A1 (n_0_2_18), .A2 (\accumulator[8] ), .B1 (n_0_9), .B2 (sps__n13));
OAI22_X1 i_0_2_52 (.ZN (n_0_332), .A1 (n_0_2_20), .A2 (n_0_2_33), .B1 (n_0_2_21), .B2 (n_0_2_34));
INV_X1 i_0_2_51 (.ZN (n_0_2_34), .A (n_0_134));
INV_X1 i_0_2_50 (.ZN (n_0_396), .A (n_0_2_33));
AOI22_X1 i_0_2_49 (.ZN (n_0_2_33), .A1 (n_0_2_18), .A2 (\accumulator[7] ), .B1 (n_0_8), .B2 (sps__n13));
OAI22_X1 i_0_2_48 (.ZN (n_0_331), .A1 (n_0_2_20), .A2 (n_0_2_31), .B1 (n_0_2_21), .B2 (n_0_2_32));
INV_X1 i_0_2_47 (.ZN (n_0_2_32), .A (n_0_133));
INV_X1 i_0_2_46 (.ZN (n_0_395), .A (n_0_2_31));
AOI22_X1 i_0_2_45 (.ZN (n_0_2_31), .A1 (n_0_2_18), .A2 (\accumulator[6] ), .B1 (n_0_7), .B2 (sps__n13));
OAI22_X1 i_0_2_44 (.ZN (n_0_330), .A1 (n_0_2_20), .A2 (n_0_2_29), .B1 (n_0_2_21), .B2 (n_0_2_30));
INV_X1 i_0_2_43 (.ZN (n_0_2_30), .A (n_0_132));
INV_X1 i_0_2_42 (.ZN (n_0_394), .A (n_0_2_29));
AOI22_X1 i_0_2_41 (.ZN (n_0_2_29), .A1 (n_0_2_18), .A2 (\accumulator[5] ), .B1 (n_0_6), .B2 (sps__n13));
OAI22_X1 i_0_2_40 (.ZN (n_0_329), .A1 (n_0_2_20), .A2 (n_0_2_27), .B1 (n_0_2_21), .B2 (n_0_2_28));
INV_X1 i_0_2_39 (.ZN (n_0_2_28), .A (n_0_131));
INV_X1 i_0_2_38 (.ZN (n_0_393), .A (n_0_2_27));
AOI22_X1 i_0_2_37 (.ZN (n_0_2_27), .A1 (n_0_2_18), .A2 (\accumulator[4] ), .B1 (n_0_5), .B2 (sps__n13));
OAI22_X1 i_0_2_36 (.ZN (n_0_328), .A1 (n_0_2_20), .A2 (n_0_2_25), .B1 (n_0_2_21), .B2 (n_0_2_26));
INV_X1 i_0_2_35 (.ZN (n_0_2_26), .A (n_0_130));
INV_X1 i_0_2_34 (.ZN (n_0_392), .A (n_0_2_25));
AOI22_X1 i_0_2_33 (.ZN (n_0_2_25), .A1 (n_0_2_18), .A2 (\accumulator[3] ), .B1 (n_0_4), .B2 (sps__n13));
OAI22_X1 i_0_2_32 (.ZN (n_0_327), .A1 (n_0_2_20), .A2 (n_0_2_23), .B1 (n_0_2_21), .B2 (n_0_2_24));
INV_X1 i_0_2_31 (.ZN (n_0_2_24), .A (n_0_129));
INV_X1 i_0_2_30 (.ZN (n_0_391), .A (n_0_2_23));
AOI22_X1 i_0_2_29 (.ZN (n_0_2_23), .A1 (n_0_2_18), .A2 (\accumulator[2] ), .B1 (n_0_3), .B2 (sps__n13));
OAI22_X1 i_0_2_28 (.ZN (n_0_326), .A1 (n_0_2_20), .A2 (n_0_2_19), .B1 (n_0_2_21), .B2 (n_0_2_22));
INV_X1 i_0_2_27 (.ZN (n_0_2_22), .A (n_0_128));
INV_X4 i_0_2_26 (.ZN (spt__n28), .A (n_0_2_16));
INV_X4 i_0_2_25 (.ZN (n_0_2_20), .A (n_0_453));
INV_X1 i_0_2_24 (.ZN (n_0_390), .A (n_0_2_19));
AOI22_X1 i_0_2_23 (.ZN (n_0_2_19), .A1 (n_0_2_18), .A2 (\accumulator[1] ), .B1 (n_0_2), .B2 (sps__n13));
INV_X4 i_0_2_22 (.ZN (n_0_2_18), .A (sps__n13));
INV_X1 i_0_2_21 (.ZN (n_0_325), .A (n_0_2_17));
AOI22_X1 i_0_2_20 (.ZN (n_0_2_17), .A1 (n_0_2_16), .A2 (n_0_127), .B1 (n_0_453), .B2 (\accumulator[0] ));
NOR2_X1 i_0_2_19 (.ZN (n_0_2_16), .A1 (n_0_2_15), .A2 (set_signal));
AND2_X2 i_0_2_18 (.ZN (n_0_453), .A1 (n_0_2_15), .A2 (n_0_2_8));
NOR4_X1 i_0_2_17 (.ZN (n_0_2_15), .A1 (n_0_2_12), .A2 (n_0_2_14), .A3 (spc__n22), .A4 (sps__n10));
NAND2_X1 i_0_2_16 (.ZN (spt__n25), .A1 (n_0_2_13), .A2 (\counter[5] ));
INV_X4 i_0_2_15 (.ZN (n_0_2_13), .A (spc__n16));
INV_X4 i_0_2_14 (.ZN (n_0_2_12), .A (n_0_2_11));
NOR2_X1 i_0_2_13 (.ZN (n_0_2_11), .A1 (sps__n4), .A2 (sps__n7));
AOI221_X1 i_0_2_12 (.ZN (n_0_324), .A (set_signal), .B1 (n_0_2_3), .B2 (\counter[5] )
    , .C1 (n_0_2_9), .C2 (n_0_2_10));
INV_X1 i_0_2_11 (.ZN (n_0_2_10), .A (\counter[5] ));
INV_X1 i_0_2_10 (.ZN (n_0_2_9), .A (n_0_2_3));
AND2_X1 i_0_2_9 (.ZN (n_0_259), .A1 (n_0_2_8), .A2 (n_0_2_7));
AND2_X1 i_0_2_8 (.ZN (n_0_258), .A1 (n_0_2_8), .A2 (n_0_2_6));
AND2_X1 i_0_2_7 (.ZN (n_0_257), .A1 (n_0_2_8), .A2 (n_0_2_5));
AND2_X1 i_0_2_6 (.ZN (n_0_256), .A1 (n_0_2_8), .A2 (n_0_2_4));
INV_X1 i_0_2_5 (.ZN (n_0_2_8), .A (set_signal));
NOR2_X1 i_0_2_4 (.ZN (n_0_255), .A1 (set_signal), .A2 (sps__n10));
HA_X1 i_0_2_3 (.CO (n_0_2_3), .S (n_0_2_7), .A (spc__n16), .B (n_0_2_2));
HA_X1 i_0_2_2 (.CO (n_0_2_2), .S (n_0_2_6), .A (spc__n22), .B (n_0_2_1));
HA_X1 i_0_2_1 (.CO (n_0_2_1), .S (n_0_2_5), .A (sps__n4), .B (n_0_2_0));
HA_X1 i_0_2_0 (.CO (n_0_2_0), .S (n_0_2_4), .A (sps__n7), .B (sps__n10));
AND2_X1 i_0_0_62 (.ZN (n_0_254), .A1 (\multiplier_reg[31] ), .A2 (n_0_95));
MUX2_X1 i_0_0_61 (.Z (n_0_253), .A (\multiplier_reg[30] ), .B (n_0_94), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_60 (.Z (n_0_252), .A (\multiplier_reg[29] ), .B (n_0_93), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_59 (.Z (n_0_251), .A (\multiplier_reg[28] ), .B (n_0_92), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_58 (.Z (n_0_250), .A (\multiplier_reg[27] ), .B (n_0_91), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_57 (.Z (n_0_249), .A (\multiplier_reg[26] ), .B (n_0_90), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_56 (.Z (n_0_248), .A (\multiplier_reg[25] ), .B (n_0_89), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_55 (.Z (n_0_247), .A (\multiplier_reg[24] ), .B (n_0_88), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_54 (.Z (n_0_246), .A (\multiplier_reg[23] ), .B (n_0_87), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_53 (.Z (n_0_245), .A (\multiplier_reg[22] ), .B (n_0_86), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_52 (.Z (n_0_244), .A (\multiplier_reg[21] ), .B (n_0_85), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_51 (.Z (n_0_243), .A (\multiplier_reg[20] ), .B (n_0_84), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_50 (.Z (n_0_242), .A (\multiplier_reg[19] ), .B (n_0_83), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_49 (.Z (n_0_241), .A (\multiplier_reg[18] ), .B (n_0_82), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_48 (.Z (n_0_240), .A (\multiplier_reg[17] ), .B (n_0_81), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_47 (.Z (n_0_239), .A (\multiplier_reg[16] ), .B (n_0_80), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_46 (.Z (n_0_238), .A (\multiplier_reg[15] ), .B (n_0_79), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_45 (.Z (n_0_237), .A (\multiplier_reg[14] ), .B (n_0_78), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_44 (.Z (n_0_236), .A (\multiplier_reg[13] ), .B (n_0_77), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_43 (.Z (n_0_235), .A (\multiplier_reg[12] ), .B (n_0_76), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_42 (.Z (n_0_234), .A (\multiplier_reg[11] ), .B (n_0_75), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_41 (.Z (n_0_233), .A (\multiplier_reg[10] ), .B (n_0_74), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_40 (.Z (n_0_232), .A (\multiplier_reg[9] ), .B (n_0_73), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_39 (.Z (n_0_231), .A (\multiplier_reg[8] ), .B (n_0_72), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_38 (.Z (n_0_230), .A (\multiplier_reg[7] ), .B (n_0_71), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_37 (.Z (n_0_229), .A (\multiplier_reg[6] ), .B (n_0_70), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_36 (.Z (n_0_227), .A (\multiplier_reg[5] ), .B (n_0_69), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_35 (.Z (n_0_226), .A (\multiplier_reg[4] ), .B (n_0_68), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_34 (.Z (n_0_225), .A (\multiplier_reg[3] ), .B (n_0_67), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_33 (.Z (n_0_224), .A (\multiplier_reg[2] ), .B (n_0_66), .S (\multiplier_reg[31] ));
MUX2_X1 i_0_0_32 (.Z (n_0_223), .A (\multiplier_reg[1] ), .B (n_0_65), .S (\multiplier_reg[31] ));
AND2_X1 i_0_0_31 (.ZN (n_0_222), .A1 (\multiplicand_reg[31] ), .A2 (n_0_126));
MUX2_X1 i_0_0_30 (.Z (n_0_221), .A (\multiplicand_reg[30] ), .B (n_0_125), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_29 (.Z (n_0_220), .A (\multiplicand_reg[29] ), .B (n_0_124), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_28 (.Z (n_0_219), .A (\multiplicand_reg[28] ), .B (n_0_123), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_27 (.Z (n_0_218), .A (\multiplicand_reg[27] ), .B (n_0_122), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_26 (.Z (n_0_217), .A (\multiplicand_reg[26] ), .B (n_0_121), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_25 (.Z (n_0_216), .A (\multiplicand_reg[25] ), .B (n_0_120), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_24 (.Z (n_0_215), .A (\multiplicand_reg[24] ), .B (n_0_119), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_23 (.Z (n_0_214), .A (\multiplicand_reg[23] ), .B (n_0_118), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_22 (.Z (n_0_213), .A (\multiplicand_reg[22] ), .B (n_0_117), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_21 (.Z (n_0_212), .A (\multiplicand_reg[21] ), .B (n_0_116), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_20 (.Z (n_0_211), .A (\multiplicand_reg[20] ), .B (n_0_115), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_19 (.Z (n_0_210), .A (\multiplicand_reg[19] ), .B (n_0_114), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_18 (.Z (n_0_209), .A (\multiplicand_reg[18] ), .B (n_0_113), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_17 (.Z (n_0_208), .A (\multiplicand_reg[17] ), .B (n_0_112), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_16 (.Z (n_0_207), .A (\multiplicand_reg[16] ), .B (n_0_111), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_15 (.Z (n_0_206), .A (\multiplicand_reg[15] ), .B (n_0_110), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_14 (.Z (n_0_205), .A (\multiplicand_reg[14] ), .B (n_0_109), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_13 (.Z (n_0_204), .A (\multiplicand_reg[13] ), .B (n_0_108), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_12 (.Z (n_0_203), .A (\multiplicand_reg[12] ), .B (n_0_107), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_11 (.Z (n_0_202), .A (\multiplicand_reg[11] ), .B (n_0_106), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_10 (.Z (n_0_201), .A (\multiplicand_reg[10] ), .B (n_0_105), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_9 (.Z (n_0_200), .A (\multiplicand_reg[9] ), .B (n_0_104), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_8 (.Z (n_0_199), .A (\multiplicand_reg[8] ), .B (n_0_103), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_7 (.Z (n_0_198), .A (\multiplicand_reg[7] ), .B (n_0_102), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_6 (.Z (n_0_197), .A (\multiplicand_reg[6] ), .B (n_0_101), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_5 (.Z (n_0_196), .A (\multiplicand_reg[5] ), .B (n_0_100), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_4 (.Z (n_0_195), .A (\multiplicand_reg[4] ), .B (n_0_99), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_3 (.Z (n_0_194), .A (\multiplicand_reg[3] ), .B (n_0_98), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_2 (.Z (n_0_193), .A (\multiplicand_reg[2] ), .B (n_0_97), .S (\multiplicand_reg[31] ));
MUX2_X1 i_0_0_1 (.Z (n_0_192), .A (\multiplicand_reg[1] ), .B (n_0_96), .S (\multiplicand_reg[31] ));
XOR2_X1 i_0_0_0 (.Z (n_0_191), .A (\multiplier_reg[31] ), .B (\multiplicand_reg[31] ));
datapath__0_15 i_0_14 (.p_1 ({n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, 
    n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, 
    n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, n_0_169, n_0_168, n_0_167, 
    n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161, n_0_160, n_0_159, n_0_158, 
    n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, 
    n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, 
    n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, 
    n_0_130, n_0_129, n_0_128, n_0_127}), .accumulator ({\accumulator[63] , \accumulator[62] , 
    \accumulator[61] , \accumulator[60] , \accumulator[59] , \accumulator[58] , \accumulator[57] , 
    \accumulator[56] , \accumulator[55] , \accumulator[54] , \accumulator[53] , \accumulator[52] , 
    \accumulator[51] , \accumulator[50] , \accumulator[49] , \accumulator[48] , \accumulator[47] , 
    \accumulator[46] , \accumulator[45] , \accumulator[44] , \accumulator[43] , \accumulator[42] , 
    \accumulator[41] , \accumulator[40] , \accumulator[39] , \accumulator[38] , \accumulator[37] , 
    \accumulator[36] , \accumulator[35] , \accumulator[34] , \accumulator[33] , \accumulator[32] , 
    \accumulator[31] , \accumulator[30] , \accumulator[29] , \accumulator[28] , \accumulator[27] , 
    \accumulator[26] , \accumulator[25] , \accumulator[24] , \accumulator[23] , \accumulator[22] , 
    \accumulator[21] , \accumulator[20] , \accumulator[19] , \accumulator[18] , \accumulator[17] , 
    \accumulator[16] , \accumulator[15] , \accumulator[14] , \accumulator[13] , \accumulator[12] , 
    \accumulator[11] , \accumulator[10] , \accumulator[9] , \accumulator[8] , \accumulator[7] , 
    \accumulator[6] , \accumulator[5] , \accumulator[4] , \accumulator[3] , \accumulator[2] , 
    \accumulator[1] , spw__n123}), .p_0 ({n_0_323, n_0_322, n_0_321, n_0_320, n_0_319, 
    n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, n_0_310, 
    n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, n_0_303, n_0_302, n_0_301, 
    n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, n_0_294, n_0_293, n_0_292, 
    n_0_291, n_0_290, n_0_289, n_0_288, n_0_287, n_0_286, n_0_285, n_0_284, n_0_283, 
    n_0_282, n_0_281, n_0_280, n_0_279, n_0_278, n_0_277, n_0_276, n_0_275, n_0_274, 
    n_0_273, n_0_272, n_0_271, n_0_270, n_0_269, n_0_268, n_0_267, n_0_266, n_0_265, 
    n_0_264, n_0_263, n_0_262, n_0_261, n_0_260}));
datapath__0_12 i_0_11 (.p_0 ({n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, 
    n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
    n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, 
    n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, uc_2}), .multiplicand_reg ({
    \multiplicand_reg[31] , \multiplicand_reg[30] , \multiplicand_reg[29] , \multiplicand_reg[28] , 
    \multiplicand_reg[27] , \multiplicand_reg[26] , \multiplicand_reg[25] , \multiplicand_reg[24] , 
    \multiplicand_reg[23] , \multiplicand_reg[22] , \multiplicand_reg[21] , \multiplicand_reg[20] , 
    \multiplicand_reg[19] , \multiplicand_reg[18] , \multiplicand_reg[17] , \multiplicand_reg[16] , 
    \multiplicand_reg[15] , \multiplicand_reg[14] , \multiplicand_reg[13] , \multiplicand_reg[12] , 
    \multiplicand_reg[11] , \multiplicand_reg[10] , \multiplicand_reg[9] , \multiplicand_reg[8] , 
    \multiplicand_reg[7] , \multiplicand_reg[6] , \multiplicand_reg[5] , \multiplicand_reg[4] , 
    \multiplicand_reg[3] , \multiplicand_reg[2] , \multiplicand_reg[1] , \multiplicand_reg[0] }));
datapath__0_3 i_0_3 (.p_0 ({n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
    n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 
    n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
    n_0_68, n_0_67, n_0_66, n_0_65, uc_1}), .multiplier_reg ({\multiplier_reg[31] , 
    \multiplier_reg[30] , \multiplier_reg[29] , \multiplier_reg[28] , \multiplier_reg[27] , 
    \multiplier_reg[26] , \multiplier_reg[25] , \multiplier_reg[24] , \multiplier_reg[23] , 
    \multiplier_reg[22] , \multiplier_reg[21] , \multiplier_reg[20] , \multiplier_reg[19] , 
    \multiplier_reg[18] , \multiplier_reg[17] , \multiplier_reg[16] , \multiplier_reg[15] , 
    \multiplier_reg[14] , \multiplier_reg[13] , \multiplier_reg[12] , \multiplier_reg[11] , 
    \multiplier_reg[10] , \multiplier_reg[9] , \multiplier_reg[8] , \multiplier_reg[7] , 
    \multiplier_reg[6] , \multiplier_reg[5] , \multiplier_reg[4] , \multiplier_reg[3] , 
    \multiplier_reg[2] , \multiplier_reg[1] , \multiplier_reg[0] }));
datapath i_0_1 (.p_0 ({n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, 
    n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, 
    n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, 
    n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, 
    n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
    n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, 
    n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, uc_0}), .accumulator ({\accumulator[63] , 
    \accumulator[62] , \accumulator[61] , \accumulator[60] , \accumulator[59] , \accumulator[58] , 
    \accumulator[57] , \accumulator[56] , \accumulator[55] , \accumulator[54] , \accumulator[53] , 
    \accumulator[52] , \accumulator[51] , \accumulator[50] , \accumulator[49] , \accumulator[48] , 
    \accumulator[47] , \accumulator[46] , \accumulator[45] , \accumulator[44] , \accumulator[43] , 
    \accumulator[42] , \accumulator[41] , \accumulator[40] , \accumulator[39] , \accumulator[38] , 
    \accumulator[37] , \accumulator[36] , \accumulator[35] , \accumulator[34] , \accumulator[33] , 
    \accumulator[32] , \accumulator[31] , \accumulator[30] , \accumulator[29] , \accumulator[28] , 
    \accumulator[27] , \accumulator[26] , \accumulator[25] , \accumulator[24] , \accumulator[23] , 
    \accumulator[22] , \accumulator[21] , \accumulator[20] , \accumulator[19] , \accumulator[18] , 
    \accumulator[17] , \accumulator[16] , \accumulator[15] , \accumulator[14] , \accumulator[13] , 
    \accumulator[12] , \accumulator[11] , \accumulator[10] , \accumulator[9] , \accumulator[8] , 
    \accumulator[7] , \accumulator[6] , \accumulator[5] , \accumulator[4] , \accumulator[3] , 
    \accumulator[2] , \accumulator[1] , spw__n124}), .accumulator_0_PP_0 (spw__n125)
    , .accumulator_1_PP_0 (\accumulator[1] ));
DFF_X1 \outmultiplier_reg_reg[0]  (.Q (\outmultiplier_reg[0] ), .CK (n_0_1), .D (spw__n124));
DFF_X1 \outmultiplier_reg_reg[1]  (.Q (\outmultiplier_reg[1] ), .CK (n_0_1), .D (n_0_390));
DFF_X1 \outmultiplier_reg_reg[2]  (.Q (\outmultiplier_reg[2] ), .CK (n_0_1), .D (n_0_391));
DFF_X1 \outmultiplier_reg_reg[3]  (.Q (\outmultiplier_reg[3] ), .CK (n_0_1), .D (n_0_392));
DFF_X1 \outmultiplier_reg_reg[4]  (.Q (\outmultiplier_reg[4] ), .CK (n_0_1), .D (n_0_393));
DFF_X1 \outmultiplier_reg_reg[5]  (.Q (\outmultiplier_reg[5] ), .CK (n_0_1), .D (n_0_394));
DFF_X1 \outmultiplier_reg_reg[6]  (.Q (\outmultiplier_reg[6] ), .CK (n_0_1), .D (n_0_395));
DFF_X1 \outmultiplier_reg_reg[7]  (.Q (\outmultiplier_reg[7] ), .CK (n_0_1), .D (n_0_396));
DFF_X1 \outmultiplier_reg_reg[8]  (.Q (\outmultiplier_reg[8] ), .CK (n_0_1), .D (n_0_397));
DFF_X1 \outmultiplier_reg_reg[9]  (.Q (\outmultiplier_reg[9] ), .CK (n_0_1), .D (n_0_398));
DFF_X1 \outmultiplier_reg_reg[10]  (.Q (\outmultiplier_reg[10] ), .CK (n_0_1), .D (n_0_399));
DFF_X1 \outmultiplier_reg_reg[11]  (.Q (\outmultiplier_reg[11] ), .CK (n_0_1), .D (n_0_400));
DFF_X1 \outmultiplier_reg_reg[12]  (.Q (\outmultiplier_reg[12] ), .CK (n_0_1), .D (n_0_401));
DFF_X1 \outmultiplier_reg_reg[13]  (.Q (\outmultiplier_reg[13] ), .CK (n_0_1), .D (n_0_402));
DFF_X1 \outmultiplier_reg_reg[14]  (.Q (\outmultiplier_reg[14] ), .CK (n_0_1), .D (n_0_403));
DFF_X1 \outmultiplier_reg_reg[15]  (.Q (\outmultiplier_reg[15] ), .CK (n_0_1), .D (n_0_404));
DFF_X1 \outmultiplier_reg_reg[16]  (.Q (\outmultiplier_reg[16] ), .CK (n_0_1), .D (n_0_405));
DFF_X1 \outmultiplier_reg_reg[17]  (.Q (\outmultiplier_reg[17] ), .CK (n_0_1), .D (n_0_406));
DFF_X1 \outmultiplier_reg_reg[18]  (.Q (\outmultiplier_reg[18] ), .CK (n_0_1), .D (n_0_407));
DFF_X1 \outmultiplier_reg_reg[19]  (.Q (\outmultiplier_reg[19] ), .CK (n_0_1), .D (n_0_408));
DFF_X1 \outmultiplier_reg_reg[20]  (.Q (\outmultiplier_reg[20] ), .CK (n_0_1), .D (n_0_409));
DFF_X1 \outmultiplier_reg_reg[21]  (.Q (\outmultiplier_reg[21] ), .CK (n_0_1), .D (n_0_410));
DFF_X1 \outmultiplier_reg_reg[22]  (.Q (\outmultiplier_reg[22] ), .CK (n_0_1), .D (n_0_411));
DFF_X1 \outmultiplier_reg_reg[23]  (.Q (\outmultiplier_reg[23] ), .CK (n_0_1), .D (n_0_412));
DFF_X1 \outmultiplier_reg_reg[24]  (.Q (\outmultiplier_reg[24] ), .CK (n_0_1), .D (n_0_413));
DFF_X1 \outmultiplier_reg_reg[25]  (.Q (\outmultiplier_reg[25] ), .CK (n_0_1), .D (n_0_414));
DFF_X1 \outmultiplier_reg_reg[26]  (.Q (\outmultiplier_reg[26] ), .CK (n_0_1), .D (n_0_415));
DFF_X1 \outmultiplier_reg_reg[27]  (.Q (\outmultiplier_reg[27] ), .CK (n_0_1), .D (n_0_416));
DFF_X1 \outmultiplier_reg_reg[28]  (.Q (\outmultiplier_reg[28] ), .CK (n_0_1), .D (n_0_417));
DFF_X1 \outmultiplier_reg_reg[29]  (.Q (\outmultiplier_reg[29] ), .CK (n_0_1), .D (n_0_418));
DFF_X1 \outmultiplier_reg_reg[30]  (.Q (\outmultiplier_reg[30] ), .CK (n_0_1), .D (n_0_419));
DFF_X1 \outmultiplier_reg_reg[31]  (.Q (\outmultiplier_reg[31] ), .CK (n_0_1), .D (n_0_420));
registerNbits outmultiplicand (.out ({product[31], product[30], product[29], product[28], 
    product[27], product[26], product[25], product[24], product[23], product[22], 
    product[21], product[20], product[19], product[18], product[17], product[16], 
    product[15], product[14], product[13], product[12], product[11], product[10], 
    product[9], product[8], product[7], product[6], product[5], product[4], product[3], 
    product[2], product[1], product[0]}), .clk (clk), .en (en), .inp ({\outmultiplier_reg[31] , 
    \outmultiplier_reg[30] , \outmultiplier_reg[29] , \outmultiplier_reg[28] , \outmultiplier_reg[27] , 
    \outmultiplier_reg[26] , \outmultiplier_reg[25] , \outmultiplier_reg[24] , \outmultiplier_reg[23] , 
    \outmultiplier_reg[22] , \outmultiplier_reg[21] , \outmultiplier_reg[20] , \outmultiplier_reg[19] , 
    \outmultiplier_reg[18] , \outmultiplier_reg[17] , \outmultiplier_reg[16] , \outmultiplier_reg[15] , 
    \outmultiplier_reg[14] , \outmultiplier_reg[13] , \outmultiplier_reg[12] , \outmultiplier_reg[11] , 
    \outmultiplier_reg[10] , \outmultiplier_reg[9] , \outmultiplier_reg[8] , \outmultiplier_reg[7] , 
    \outmultiplier_reg[6] , \outmultiplier_reg[5] , \outmultiplier_reg[4] , \outmultiplier_reg[3] , 
    \outmultiplier_reg[2] , \outmultiplier_reg[1] , \outmultiplier_reg[0] }), .reset (reset));
registerNbits__0_28 outmultiplier (.out ({product[63], product[62], product[61], 
    product[60], product[59], product[58], product[57], product[56], product[55], 
    product[54], product[53], product[52], product[51], product[50], product[49], 
    product[48], product[47], product[46], product[45], product[44], product[43], 
    product[42], product[41], product[40], product[39], product[38], product[37], 
    product[36], product[35], product[34], product[33], product[32]}), .clk (clk)
    , .en (en), .inp ({\outmultiplicand_reg[31] , \outmultiplicand_reg[30] , \outmultiplicand_reg[29] , 
    \outmultiplicand_reg[28] , \outmultiplicand_reg[27] , \outmultiplicand_reg[26] , 
    \outmultiplicand_reg[25] , \outmultiplicand_reg[24] , \outmultiplicand_reg[23] , 
    \outmultiplicand_reg[22] , \outmultiplicand_reg[21] , \outmultiplicand_reg[20] , 
    \outmultiplicand_reg[19] , \outmultiplicand_reg[18] , \outmultiplicand_reg[17] , 
    \outmultiplicand_reg[16] , \outmultiplicand_reg[15] , \outmultiplicand_reg[14] , 
    \outmultiplicand_reg[13] , \outmultiplicand_reg[12] , \outmultiplicand_reg[11] , 
    \outmultiplicand_reg[10] , \outmultiplicand_reg[9] , \outmultiplicand_reg[8] , 
    \outmultiplicand_reg[7] , \outmultiplicand_reg[6] , \outmultiplicand_reg[5] , 
    \outmultiplicand_reg[4] , \outmultiplicand_reg[3] , \outmultiplicand_reg[2] , 
    \outmultiplicand_reg[1] , \outmultiplicand_reg[0] }), .reset (reset));
registerNbits__0_25 regmultiplier (.out ({\multiplier_reg[31] , \multiplier_reg[30] , 
    \multiplier_reg[29] , \multiplier_reg[28] , \multiplier_reg[27] , \multiplier_reg[26] , 
    \multiplier_reg[25] , \multiplier_reg[24] , \multiplier_reg[23] , \multiplier_reg[22] , 
    \multiplier_reg[21] , \multiplier_reg[20] , \multiplier_reg[19] , \multiplier_reg[18] , 
    \multiplier_reg[17] , \multiplier_reg[16] , \multiplier_reg[15] , \multiplier_reg[14] , 
    \multiplier_reg[13] , \multiplier_reg[12] , \multiplier_reg[11] , \multiplier_reg[10] , 
    \multiplier_reg[9] , \multiplier_reg[8] , \multiplier_reg[7] , \multiplier_reg[6] , 
    \multiplier_reg[5] , \multiplier_reg[4] , \multiplier_reg[3] , \multiplier_reg[2] , 
    \multiplier_reg[1] , \multiplier_reg[0] }), .clk (clk), .en (en), .inp ({multiplier[31], 
    multiplier[30], multiplier[29], multiplier[28], multiplier[27], multiplier[26], 
    multiplier[25], multiplier[24], multiplier[23], multiplier[22], multiplier[21], 
    multiplier[20], multiplier[19], multiplier[18], multiplier[17], multiplier[16], 
    multiplier[15], multiplier[14], multiplier[13], multiplier[12], multiplier[11], 
    multiplier[10], multiplier[9], multiplier[8], multiplier[7], multiplier[6], multiplier[5], 
    multiplier[4], multiplier[3], multiplier[2], multiplier[1], multiplier[0]}), .reset (reset));
registerNbits__0_22 regmultiplicand (.out ({\multiplicand_reg[31] , \multiplicand_reg[30] , 
    \multiplicand_reg[29] , \multiplicand_reg[28] , \multiplicand_reg[27] , \multiplicand_reg[26] , 
    \multiplicand_reg[25] , \multiplicand_reg[24] , \multiplicand_reg[23] , \multiplicand_reg[22] , 
    \multiplicand_reg[21] , \multiplicand_reg[20] , \multiplicand_reg[19] , \multiplicand_reg[18] , 
    \multiplicand_reg[17] , \multiplicand_reg[16] , \multiplicand_reg[15] , \multiplicand_reg[14] , 
    \multiplicand_reg[13] , \multiplicand_reg[12] , \multiplicand_reg[11] , \multiplicand_reg[10] , 
    \multiplicand_reg[9] , \multiplicand_reg[8] , \multiplicand_reg[7] , \multiplicand_reg[6] , 
    \multiplicand_reg[5] , \multiplicand_reg[4] , \multiplicand_reg[3] , \multiplicand_reg[2] , 
    \multiplicand_reg[1] , \multiplicand_reg[0] }), .clk (clk), .en (en), .inp ({
    multipicand[31], multipicand[30], multipicand[29], multipicand[28], multipicand[27], 
    multipicand[26], multipicand[25], multipicand[24], multipicand[23], multipicand[22], 
    multipicand[21], multipicand[20], multipicand[19], multipicand[18], multipicand[17], 
    multipicand[16], multipicand[15], multipicand[14], multipicand[13], multipicand[12], 
    multipicand[11], multipicand[10], multipicand[9], multipicand[8], multipicand[7], 
    multipicand[6], multipicand[5], multipicand[4], multipicand[3], multipicand[2], 
    multipicand[1], multipicand[0]}), .reset (reset));
BUF_X8 sps__L1_c1 (.Z (sps__n1), .A (n_0_2_149));
BUF_X8 sps__L1_c4 (.Z (sps__n4), .A (\counter[2] ));
BUF_X8 sps__L1_c7 (.Z (sps__n7), .A (\counter[1] ));
BUF_X8 sps__L1_c10 (.Z (sps__n10), .A (\counter[0] ));
BUF_X8 sps__L1_c13 (.Z (sps__n13), .A (negative_product_flag));
BUF_X8 spc__L1_c16 (.Z (spc__n16), .A (\counter[4] ));
BUF_X8 spc__L1_c19 (.Z (spc__n19), .A (n_0_2_147));
BUF_X8 spc__L1_c22 (.Z (spc__n22), .A (\counter[3] ));
BUF_X4 spt__c25 (.Z (n_0_2_14), .A (spt__n25));
BUF_X16 spt__c28 (.Z (n_0_2_21), .A (spt__n28));
CLKBUF_X1 spw__L2_c2_c123 (.Z (\accumulator[0] ), .A (spw__n123));
CLKBUF_X1 spw__L1_c1_c124 (.Z (spw__n123), .A (spw__n125));
CLKBUF_X1 spw__L1_c4_c125 (.Z (spw__n124), .A (spw__n125));
BUF_X2 spw__L1_c155 (.Z (spw__n155), .A (sps__n1));
CLKBUF_X3 spw__L2_c156 (.Z (spw__n156), .A (spw__n155));
BUF_X1 spw__L1_c325 (.Z (spw__n309), .A (sps__n7));
BUF_X2 spw__L2_c326 (.Z (spw__n310), .A (spw__n309));
BUF_X2 spw__L3_c327 (.Z (spw__n311), .A (spw__n310));
BUF_X2 spw__L2_c328 (.Z (spw__n312), .A (spw__n309));
BUF_X2 spw__L1_c339 (.Z (spw__n323), .A (n_0_2_148));
BUF_X2 spw__L1_c340 (.Z (spw__n324), .A (n_0_2_148));
CLKBUF_X3 spw__L2_c341 (.Z (spw__n325), .A (spw__n324));
BUF_X2 spw__L3_c342 (.Z (spw__n326), .A (spw__n325));
BUF_X2 spw__L1_c353 (.Z (spw__n337), .A (sps__n4));
CLKBUF_X3 spw__L2_c354 (.Z (spw__n338), .A (spw__n337));

endmodule //sequential_multiplier


